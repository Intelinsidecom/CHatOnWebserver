.                                                                                                                                    	                                                      	   	                                 -       	                                                                                                                                                                                                    -                                                                                                                                                                                                                                  ,                                                                                                                                    
	                                                                                 2                               	                                                       	                                                                                                                              .                                                                                                                                                                                                            	                -                                                                                                                                                                                                                2               	                                                                                                                                                                                                /                                                                                                                                   	                                                                                   -                                                                                                                                                                                                           	          /                                                                                                                                                                                                    
       /                                                                                                                                                                                                                   2                                                                                                                                                                                                               .                                                                                                                                                                                                             -                                                                                                                                                                                                                
       
  -                                                                                                                                                                                                                    ,                                                                                                                                                                                                                              -                                                                                        	 
                                                                                                                                        ,              	                                                                                                                     	                                                                                         ,                                                                                                                                                                                                               /                                                                                                                                                                                                                        ,                                                                                                                                                                                                                         
   -                                                                                                                                                                                                        /                                                                                                                                                                                                                         0                                                                                                                                                                                                                     	.          
                                                                                                                                                                                                        .                                                                                                                                                                                                             .   
                                                                                                                                                                                                                       0                                                                                       
                                                                                                                 	.                                                                                                                                                                                                                                   -                                                                                                                                                                                                                                     0                                                                                                                              	                                                                                          1                                                                                                                                                                                                            -                                                                                                                                                                                                                    -                                                                                                                                                                                            
 
                                   1                                                                                                                                                                                                         /                                                                                                                                                                                                                /                                                                                                                                                                                                       /                                                                                                                                                                                                      0               	                                                                                                                  
                                                                                           1                                                                                                                                                                                                                
           -                                                                                                                                                                                                                   	           0                                                                                                                                                                                                     - 	                         	                                                                                                                                                                                            1                                                                                                                                                                                                     
             .                                                                                                                                                                                                                   -        	                                                                                                                                                                                                                         0                                                                                                                                                                                                          1                                                                                                                                                                                          	                            
  -                                                                                                                                                                                                                  	,                                                                                                                                                                                                                              	          -                                                                                                                                                                                                                /                                                                                    
                                                                                                                                 -       	                                                                                                                                                                                                                         ,                                                                                                                                                                                                              
                   /                                                                                                                                                                                                         ,                                                                                                                                       	                                                        
                             .               	                                                                                                                                                                                                                     /                                                                                                                                                                                                   	       
           3                                                                                                                                                                                                             	     1                                                                                                                                                                                                              .                                                                                                                                                                                                                    .                                                                                                                                                                                                             
     	          	  0                                                                                                                                                                                                                   .                                                                                                                                                                                                                          -                                                                                                                                                                                                                        ,                                                                                                                                       
                                                                                         .                                                                                                                                                                                                           ,                                                                                                                                                                                                                                 .                                                                                                                                                                                                                 	   -                                                                                                                                                                                                         -                                                                                                                                                                                                                           0                                                                                                                                                                                                                    .                                                                                                                                  	
                                                                                         0                                                                                                                                                                                                            -                                                                                                                                                                                                                                 1                                                                                                                                                                                                                 /                                                                                                                                                                                                                       0                               	                                                                                                                                                                                                .                                                                                        	                                                                                                                         3                                                                                                                                                                                                        -                                                                                                                                                                                                                   .                                                                                                                                                                                                                       2                                                                                                                                                                                                                0                                                                                                                                                                                                                .                                                                                                                                                                                                                 /                                                                                                                                                                                                   .                                                                                                                                                                                                                             .                                                                                                                                                                                                     
                    /                                                                                                                                                                                                        
              -                                                                                                                                                                                                            -                                                                                                                                                                                                                              1                	                                                                                                                                                                                                  -                                                                                                                                                                                                                                ,     
                                                                                  
                                                                                                                                              -                                                                                                                                                                                                                   /                                                                                                                                                                                        #                                 -                                                                                                                                                                                                                          .                                                                                                                                                                                                       
                   .                                                                                                                                                                                                                                ,                                  	   
                                                                                                                                                                         
               -              	                                                                                                                                                                                                                      ,                                                                                                                                                                                                                            .                                                                                                                                                                                                                           .                                                                                                                                                                                                                -                                                                                                                                                                                                              .                                                                                                                                                                                                                   	     
   .                                                                                                                                                                                                                             	  0                                                                                                                                                                                                                 .                	                                                                                                                                                                                                           -                                                                                                                                                                                                                   	1         	                                                                                                                                                                                                            -                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                /                                                                                                                                                                                                                   -                	                                                                                                                                                                                                            .                                                                                                                                                                                                                            -                                                                                                                                                                                                    	            .                                                                                                                                                                                                     
          -    
                                                                                                                                                                                                                   /                                                                                                                                                                                                                   /                                                                                                                                                                                                                               -                                                                                                                                                                                                                        -    	                                                                                                                                                                                                                        3                                                                                                                                                                                                              0                                                                                                                                                                                                               2                                                                                                                                                                                                          .                                                                                           
                                                                                                                                .                                                                                                                                                                                                               2                                                                                                                                                                                                /                                                                                                                                                             	                                                     .                                                                                                                                                                                                                      1                                                                                                                                                                                                                   /                                                                                                                                                                                                           1                                                                                                                                                                                       
                              -                                                                                                                                     
                                                                                          .                                                                                                                                                                                                                       0                                                                                                                                                                                                             	.                                                                                                                                                                                                         
           .   	                                                                                                                                                                                                                       /                                                                                                                                                                                                                     .                                                                                                                                         
                                                                          
     /                                                                                                                                                                                                                      .                   
                                                                                                                                                                                                            .                                                                                                                                                                                                                            .                                                                                                                                                                                                                    /                                                                                                                                                                                                          
        	  .            
                                                                                                                                                                                                                -                               
                                                                                                                                                                                          -        	                     
                                                                                                                                                                                              -                                                                                                                                                                                                                         0                                                                                                                                                                                                                             1                                                                                                                                                                                                           ,                                                                                                                                                                                                  
           /                                                                                                                                                                                                                       ,                                                                                                                                                                                                            
      
            .                                                                                                                                                                                                         /                                                                                                                                                                                                                        /                                                                                                                                                                                                                   	/                                                                                                                                                                                                                           -                                                                                                                                                                                                          
       -                                                                                                                                                                                                                             .                                                                                                                                                                                                                  .            	                                                                                                                                                                                                                  .                                                                                                                                                                                                                        .                                                                                                                                                                                                                           /                                                                                                                                                                                                              .             
                                                                                                                                                                                                             .                                                                                                                                                                                                                   /                     	                                                                                                                                                                                                     -                                                                                                                                                                                                                                ,                 	                                                                                                                                                                                                             .                                                                                                                                                                                                           .                                                                                                                                                                                                       /                                                                                                                                                                                                                   ,                                                                                                                                                                                                                           .                                                                                                                                                                                                               /                                                                                                                                                                                                        -                                                                                                                      
                                                                                         /                                                                                              	                                                                                                                     .                                                                                                                                                                                                                -                                                                                                                                                                                                       .                                                                                                                                                                                                                           -                                                                                                                                        
                                                                                                 /                                                                                                                                                                                                        	    
        /                                                                                                                                                                                                      
.                                                                                                                                                                                                                 /            	       	                                                                                                                                                                                                     -                                                                                                                                                                                                                       /                                                                                                                                                                                                                   	        -                                                                                                                                                                                                                            ,                                                                                                                                                                                                                       -                                                                                                                                                                                                                 
        .                                                                                                                                                                                                               2                                                                                                                                                                                                                 	.           $                                                                                                                                                                                                                        0                                                                                                                                                                                                              /           	                                                                                                                                                                                                        .                                                                                                                                                                                                                       .                                                                                                                                                                                                                             .               	                                                                                                                                                                                     .         	                                                                                                                                                                                      	               .                                                                                                                                                                                                                    /                                                                                                                                                                                                                         1                                                                                                                                                                                                 	             .      	                                                                                                                                                                                                         .                                                                                                                                                                                                              
.                                                                                                                                                                                                                     -                                                                                                                                                                                                                    -                                                                                                                                                                                                              	                -                                                                                                                                                                                    
                           .                    	                                                                                                                                                                                                        /        
                                                                                                                                                                                                            
         .                                                                                                                                                                                                                .                                                                                                                                                                                                  	            0       
       
                                                                                                                                                                                                             .                                                                                                                                                                                                                  .                                                                                                                                                                                                                                    -                                                                                             	                                                                                                                            -                            
                                                                                                                                                                                               .                                                                                                                                                                                                                  1                                                                                     	                                                                                                                      /                                                                                     	                                                                                                                              ,                                                                                                                                                                                             
                                1                                                                                                                                                                                      
                             2                                                                                                                                                                                                      0                                                                                                                                                                                                                       .                                                                                                                                                                                                             	             .                                                                                                                                                                                                     
             0                                                                                                                                                                                                   .                                                                                                                                                                                                                         .                                                                                                                                                                                                                                /                                                                                                                                                                                                               	     
   1                                                                                                                                                                                                             
.                                                                                                                                                                                                     
             .     	              	                                                                                                                                                                                                           -                                                                                                                                                                                                            /                                                                                                                                                                                                                    .                                                                                       	                                                                                                                             /                                                                                                                                                                                                                            /                                                                                                                                                                                                                    /               
                                                                                                                                                                                                       -                                                                                                                                                                                                          .                                                                                                                                                                                                                           -                                                                                                                                                                                                                        -                 	                                                                                                                                                                                                           -                                                                                                                                                                                                         .                                                                                                                                                                                                          
            .                                                                                                                                                                                                                     /         	                                                                                                                                                                                                         2                                                                                                                                                                                                             0                                                                                                                                                                                                              /                                                                                                                                                                                                    	             ,                                                                                                                                                                                                                   /                                                                                                                                                                                                         1                                                                                                                                                                                                                   -                                    :                                                                                                                                                                                                 0                                                                                                                                                                                                                         .                                                                                                                                                                                                         ,                    
                                                                                                                                                                                             0                                                                                                                                                                                                                         ,                                                                                                                                                                                                     
/                                                                                                                                                                                                           /                                                                                                                                                                                                           -                                                                                         	                                                                                                                                           -                                                                                                                                                                                                                     .                                                                                                                                                                                                  	             ,                                                                                                                                                                                                                          0                                                                                                                                                                                                                   .                                                                                                                                                                                                                               ,    	                            	                                                                                                                                                                                             /                                                                                              	                                                                                                                            4                                                                                                                                                                                                       -                                                                                                                                                                                          	                        ,                                                                                                                                                                                                                           .                                                                                                                                                                                                             	      -                                                                                                                                                                                                                            /                                                                                                                                                                                                    
.                                                                                                                                                                                                                      .                                                                                                                          
                                                                                         -         	                                                                                                                                                                                                  
                        /                                                                                                                                                                                                       0                                                                                                                                                                                                             0                	                                                                                                                                                                                                   ,                                                                                                                                                                                                                 	            -                                                                                                                                                                                                                         .                                                                                     
                                                                                                                           -                                   
                                                                                                                                                                                  .                                                                                                                                                                                                                       -                                                                                                                                                                                                                        1                                                                                                                                                                                                               .                                                                                                                                                                                                                             /                                	                                                        	                                                                                                                                  -                                                                                                                                                                                                                                   -                                                                                                                                                                                                        
    -                                                                                                                                                                                                                           -                                                                                                                                                                                                                        0                                                                                                                                                                                                                          0                                                                                                                                                                                                             .                                                                                                                                                                                                                               /                                                                                                                                                                                                 		               -                                                                                                                                                                                                                           /                                                                                                                                                                                                                    /                                                                                                                                                                                                                    -                                       9                                                            	                                                                                                                                     0                                                                                                                                                                                                                      -           	                                                                                                                                                                                                          .                                 	                                                        
                                                                                                                             /                                                                                                                                                                                                                              3                                                                                                                                                                                                              .                                                                                                                                                                                                               /          
      
                                                                                                                                                                                                 ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                           /                                                                                        	
                                                                                                                             -   	                                                                                                                                                                                                                /                                                                                    	                                                                                                                           ,                                                                                       	                                                                                                                              /                                                                                     	                                                                                                                                    /                                                                                      
                                                                                                                               /                                                                                                                                                                                                           1                                                                                                                                                                                                              
-                                                                                                                                                                                                                           	.                                                                                                                                                                                                                  .                                                                                                                                                                                                                            0                                                                                                                                                                                                  .                                                                                                                                                                                     
                                  /                                                                                                                                                                                                                      .                    	                                                                                                                                                                                                  	            /                                                                                                                                                                                                         /                                                                                                                                                                                                                0                                                                                                                                                                                                                     ,                                                                                                                                                                                                                      
             /                                                                                                                                                                                                                           -                                                                                                                                                                                                                        	    .       	                       
                                                                                                                                                                                           	.                                                                                                                                                                                                                               -                                                                                                                                                                                                                             .                                                                                                                                                                                                            -                                                                                                                                                                                                                       -                               	                                                                                                                                                                                        ,    	         	                                                                                                                                                                                                                    /                                                                                                                                                                                                        	         /                                                                                                                                                                                                                           
    /                                                                                                                                                                                                                   .             	                                                                                                                                                                                                    	           .                                                                                                                                                                                                    	         /                                                                                                                                                                                                                            /                                                                                                                                                                                                                               .                                 	                                                                                                                                                                                 	              -                                                                                                                                                                                                                     .                                                                                                                                                                                                                     ,                                     8                                                                                                                                                                                                 /    	                             	                                                                                                                                                                                        -                                                                                                                                                                             	                               .                                                                                                                                                                                                                  .                                                                                                                                                                                                                         0                                                                                                                                                                                                      
0                                                                                                                                                                                                            -  	            
                                                                                                                                                                                                     /                                                                                                                                                                                                                               /                	      	                                                                                                        	                                                                                            /                                                                                      
                                                                                                                            .     	                                                                                                                                                                                                                     /                                                                                    	                                                                                                                            -                                                                                           	                                                                                                                               1                                                                                  	                                                                                                                               /                                                                                                                                                                                     
                                1                                                                                                                                                                                                            1                                                                                                                                                                                                                

1                                                                                                                                                                                                                   .                                                                                                                                                                                                                      .                 
                                                                                                                                                                                                              /                                                                                                                                                                                                     	0                                                                                                                                                                                                                        .          
                                                                                                                                                                                                         ,        	                                                                                                                                                                                                                    /                                                                                                                                                                                               /                                                                                                                                                                                                            0    	                                                                                                                                                                                                                     ,                                                                                                                                                                                                                             0                                                                                                                                      

                                                        	                          /                                                                                                                                                                                                                       0      	   
                                                                                                                                                                                                                -                                                                                                                                                                                                                            .                                                                                                                                                                                                                     .                                                                                                                                                                                                                             "       .                                                                                                                                                                                                                   ,                                                                                                                                                                                                        	              /       	                                                                                                                                                                                                                    -                                                                                                                                                                                                                                     
    0                                                                                                                                                                                                                    .                                                                                                                                                                                                                      .                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                           .               
   
                                                                                                                                                                                                    .                   	                                                                        
                                                                                                                            .                                                                                                                                                                                                      .                                                                                                                                                                                                                     (              -       	                                                                                                                                                                                                                  0                                                                                                                                                                                                         /                                                                                                                                                                                                            -                                                                                                                                                                                                          .                                                                                                                                                                                                        0                                                                                                                                                                                                                              -                                                                                                                                                                                                                
	          0                                                                                                                                                                                                        ,                                                                                                                                                                                                                                   .                                                                                                                                                                                                          "               ,     	            
                                                                                                                                                                                                        -                                                                                                                                                                                                        /                                                                                                                                                                                                                    2                                                                                                                                                                                                 	            
-                                                                                       
                                                                                                                                0                                                                                                                                                                                        
                                 0                                                                                                                                                                                                                    0                                                                                                                                                                                                               /                                                                                                                               	                                                      
                           	-                                                                                                                                                                                        
                      .                                                                                                                                                                                                          -                                                                                                                                                                                                                    ,                                                                                                                                                                                                                  	  1                                                                                                                                    
                                                                                         ,                                                                                                                                                                                                                             0                                                                                                                                                                                                             	              -                                                                                                                                                                                                                 
        
 -                                                                                                                                                                                           
              -            
      
                                                                                                                                                                                                              1                                                                                      	                                                                                                                     /                                                                                                                                                                                        
                         -                                                                                      
                                                                                                                                    .                                                                                                                                                                                                                     /                                                                                                                                                                                                                                 .                                                                                                                                                                                                                     ,                                                                                                                                                                                                                               %      /                                                                                                                                                                                                                     .                                                                                                                                                                                                                          .         	                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                         .                                                                                                                                                                                                                             -                                                                                                                                                                                                                 -                                                                                                                                                                                                                        ,                                                                                                                                                                                                                 	              
     /   	                                                                                                                                                                                                                     /                                                                                                                                                                                                                    /                                                                                                                                                                                                                     -                                                                                                                                                                                                                    )	              /                                                                                                                                                                                                                           /                                                                                                                                                                                                 	-                                                                                                                                                                                                                 .                                                                                                                         
                                                                                         /                                                                                                                                                                                                  -                                                                                                                                                                                                                                 -                                                                                                                                                                                                               	           .                                                                                                                                                                                                         /                                                                                                                                                                                                                                 -                                                                                                                                                                                                          +                ,     	                                                                                                                                                                                                      
                 .                                	                                                                                                                                                                                -    
                                                                                                                                                                                                               0                                                                                                                                                                                                               	0                                                                                                                                                                                                                            ,                                                                                            	                                                                                                                                   1                                                                                                                                                                                                                      -                                                                                                                                                                                                        ,                                                                                                                               	                                                   	                          .                                                                                                                                                                                                                        1                                                                                                                                                                                                       .          	                                                                                                                                                                                                                    ,                                                                                                                                                                                                                          -                                                                                                                                    
                                                                                        -               
                                                                                                                                                                                                                    .                    	                                                                                                                                                                                         	                      .                                                                                                                                                                                                                                 /                                                                                                                                                                                                    -                                                                                                                                                                                                                                        /                                                                                                                                                                                                             -                                                                                                                                                                                                                        -                                                                                         
                                                                                                                                       -                                                                                                                                                                                                                .                                                                                                                                                                                                                         .                                                                                                                                                                                                                ,                                                                                                                                                                                                                               +      .            
                                                                                                                                                                                                              -                                      	                                                                                                                                                                           	             -                                 	                                                                                                                                                                                              .                                                                                                                                                                                                                                       /          	                                                                                                                                                                                          	           -          
                                                                                                                                                                                                               ,                                                                                                                                                                                                             .                                                                                                                                                                                                                                   -                                                                                                                                                                                                                                0                                                                                                                                                                                                   	             -                                                                                                                                                                                                                 ,                                                                                                                                                                                                                       1           /        #                                                                                                                                                                                                              2                                                                                                                                                                                                          ,                                                                                                                                                                                                                  .              	                                                                                                                                                                                                       1                                                                                                                                                                                                              /                                                                                                                                                                                                                                 -                                                                                                                                                                                                                           
   .                                                                                                                                                                                                    .                                                                                                                                                                                                                                    .                                                                                                                                                                                                             *                 ,                         
                                                                                                                                                                                                    /                            	                                                                                                                                                                               .        	              	                                                                                                                                                                                                  0                                                                                                                                                                                                           .                                                                                                                                                                                                                     ,                                                                                             
                                                                                                                                0                                                                                                                                                                                                                            -                                                                                                                                                                       	                            -                                                                                                                                                                                                                 	.                                                                                                                                                                                                                 .                                                                                         	                                                                                                                      /                                                                                                                                                                                                                        -                                                                                                                                                                                                                 .                                                                                                                                                                                                	                             ,   	           	                                                                                                                                                                                                            .                                                                                                                                                                                                         	                    -                                                                                                                                                                                                                	              	   0                                                                                                                                                                                                        -          	                                                                                                                                                                                                                          0                                                                                                                                                                                                             ,                                                                                                                                     	                                                                                  -       
                                                                                                                                                                                                                          /                                                                                                                                                                                                              0                                                                                                                                                                                                                            .              
                                                                                                                                                                                                  /                                                                                                                                                                                                                   
  -               
                                                                                                                                                                                                           -                                                                                         	                                                                                                                                 /       
     
                                                                                                                                                                                                               -                                                                                                                                                                                                                                   /                                                                                                                                                                                                                               ,                                                                                                                                                                                                         
     
         ,                                                                                                                                                                                                                      -                                                                                                                                                                                                                  
                   .                                                                                                                                                                                                                                   0                                                                                                                                                                                                                /      
                                                                                                                                                                                                           1                                                                                                                                                                                                                 !    	    	   ,                              	                                                                                                                                                                                       -                                                                                                                                                                                                                   -                                                                                       
 
                                                                                                                                           .                                                                                                                                                                               	                         .                                                                                                                                                                                                                  -                                                                                                                                                                                                                            /                 	                                                                                                                                                                                                  4                                   	                                                                                                                                                                          -   
          	                                                                                                                                                                                                     -                                                                                                                                                                                                                  %               ,                                                                                                                                   
                                                                                              0                                                                                                                                                                                                     ,                                                                                                                                                                                                                      .                                                                                                                                                                                                          /                                                                                                                                                                                                                          /                                                                                             	                                                                                                                            0                                                                                           
                                                                                                                                .                                                                                                                                                                                                       -                                                                                                                                                                                                 /                                                                                                                                                                                                                1                                                                                                                                                                                                  -                                                                                                                                                                                                                                0                                                                                                                                                                                                            /                                                                                                                                                                                                          -                                                                                                                                                                                                                            .                     
                                                                                                                                                                                      
                           0                                                                                                                                                                                                              .                                                                                                                                                                                                       -                                                                                                                                                                                                                        0                                                                                                                                                                                                               %             2                                                                                                                                                                                                                 /                                                                                                                                                                                                                         -                                                                                                                                                                                                               -                                                                                                                                                                                                                    -                                                                                                                                                                                                                /                                                                                                                                                                                                                           0                                                                                                                             	                                                                                           -                                                                                                                                                                                                                          -                                                                                                                                                                                                                              -                                                                                                 	                                                                                                                            	  -               	      	                                                                                                                                                                                                         .                                                                                                                                                                                                                ,                                                                                                                                                                                                                               -                                                                                                                                                                                                                
      
            .                  	                                                                                                                                                                                                                 .                                                                                                                                                                                                                              .                                                                                                                                                                                                     .                                                                                                                                                                                                            	               
  -                              
                                                                                                                                                                                            -                                                                                                                                                                                                                         -      	                                                                              	 	                                                                                                                                      /                                                                                                                                                                             
                              -                            
                                                                                             	                                                                                           /                      
                                                                                                                                                                                                             .                                                                                                                                                                                                               .                                                                                                                                                                                                             .                 
                                                                                                                                                                                                     -         
             	                                                                                                                                                                                                 !                  ,                                                                                                                                                                                                                        0                              
                                                                                                                                                                                -                                	                                                                                                                                                                                           /                                                                                                                                                                                                                         .                                                                                                                                                                                                            
            /                                 	 	                                                                                                                                                                                          /                                                                                                                                                                                                                       1                                                                                                                                                                                                      
.                                                                                                                                                                                                           0                                                                                                                                                                                    
                            0                                                                                                                                                                                                            -                                                                                                                                                                                                 	                              /            	                                                                                                                                                                                                          0                                                                                                                                                                                                            -           
                                                                                                              
                                                                                         ,                                                                                                                                                                                                                         
    -                                    	                                                                                                                                                                                 1                                                                                                                                                                                                            -                                                                                                                                                                                                                         .                                                                                                                                                                                                             
       !              -                                                                                                                                                                                                            .                                                                                  	                                                                                                                                      .                                                                                                                                                                                                                      -                                                                                                                                                                                                                   .             
                                                                                                                                                                                                       	.                                                                                                                                                                                                                     	  -                                                                                                                                                                                                                         .                                                                                                                                                                                                                     -                                                                                                                                                                                                                        .                                                                                                                                                                                                                     
      
  -                    	                                                                                                                                                                                  
                 /                                                                                                                                                                                                   	        ,                                                                                                                                                                                                                      ,                                                                                                                                                                                                                    
        -                                                                                                                                                                                                                          -              	                                                                                                                                                                                        	                0         
                                                                                                                                                                                                     .                                                                                                                                                                                                                             .                               
                                                                                                                                                                                      ,                                     
                                                                                                                                                                                    ,                                                                                   
                                                                                                                                         /                                                                                                                                                                                                          ,                    	                                                                                                                                                                                                   /         
                                                                                                                                                                                                                 -                                                                                                                                                                                                              
          0                                                                                                                        	                                                                                      0            	      
                                                                                                                                                                                                              -                                                                                                                                                                                                                        $                 ,                                                                                                                                 	                                                                                             /                                                                                                                                                                                                         ,         	                                                                                                                                                                                                                   .                                                                                                                                                                                                                         .                                                                                                                                                                                                                         -                                      
 
                                                          	                                      
                                                                                        2                                                                                                                                                                                                                    /                                                                                                                                                                                                  .                                                                                         
                                                                                                                    -                                                                                                                                                                                                                        0                                                                                                                                                                                                           ,                                                                                                                                                                                                
                          #      .                                                                                                                                                                                                               0                                                                                                                                                                                                               -                                                                                                                                 
                                                                                           /                                                                                                                                                                                                                              	       .                                                                                                                                                                                                                     2                                	                                                                                                                                                                             -                                                                                                                                                                                                                           .                                                                                                                                                                                                                   #              ,                                                                                                                                       
                                                                              .                                                                                   	                                                                                                                  
                -                            	                                                                                                  	                                                                                         ,                                                                                                                                                                                                       	                            	      ,                                                                                                                                                                                                                                 -                                       
                                                                                                                                                                              
     .                                                                                                                                                                                                                    
                          .                                                                                                                                                                                                                        
       .         
    
                                                                                                                                                                                                             .                                                                                                                                                                                                                                ,                                                                                                                                                                                                                       '         .                                                                                                                                                                                                                                -           
           	                                                                                                                                                                                              	          -                                                                                                                                                                                                                                   -                                                                                                                                                                                                                                  -                                                                                                                                                                                                                 '               ,                                                                                                                                                                                                                             -                                                                                                                                                                                                              	       -                                                                                                                                                                                                                                         .                                                                                                                                                                                                                    
          ,                                                                                                                                                                                                                                   -                                                                                                                                                                                                                               -                                                                                                                                                                                                                   -                                                                                                                                                                                                                                           ,                 1                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                             0                                                                                                                                                                                                            
,                                                                                                                                                                                                                             "             ,                                                                                         	                                                                                                                                                -                                                                                                                                                                                                                              -       
                                                                                                                                                                                                                 ,                                                                                                                                                                                                                         	                 ,                                                                                                                                                                                                                                             -            
                                                                                                                                                                                                                           -                                                                                                                                                                                                                   ,                                                                                                                                                                                                                           	         
  ,                                                                                                                                                                                                                                           -                                                                                                                                                                                                                           /                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                  "         ,             )           
                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                     .                                                                                                                                                                                                        	                 -                        
                                                                                                                                                                                                        ,                     
                                                                                                                                                                                                                    /                                                                                                                                                                                                                                   
    -                                                                                                                                                                                                     
               ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                        -                  
                                                                                                                                                                                                  	               ,                                                                                             
                                        	                                                                                        -                                                                                                                                                                                                                       
         ,                                                                                                                                                                                                                          -                                                                                                                                                                                                                                  	     ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                       (     
    ,                                                                                                                                                                                                                               .                                                                                                                                                                                                                               0                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                ,                
                                                                                                                                                                                                              .                                                                                                                                                                                                                       
               -                                                                                                 	                                                                                                                                   -                                                                                         
	                                                                                                                  
             ,                                                                                                                                                                                                                 -                                                                                                                                                                                                                             -                                                                                                                                                                                             	                            .                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                         -                                                                                                                                                                                                                               -                                                                                                                                                                                                                           %           ,                                                                                                                                                                                                                                     .            	                                                                                                                                                                                                                       -          	                                                                                                                                                                                                          ,                                                                                                                                                                                                                            7                    ,                                                                                                                                                                                                                                         ,                                                                                                                                                   
                                                                                              -                                  
                                                                                                                                                                                                      ,                                                                                                                                                                                                                                   "                ,                                                                                              	                                                                                                                        
              ,                                   :   
                                                                                                                                                                                                          ,                                                                                                                                                                                                                             
                    ,                                                                                                                                                                                                                              	         	   	     ,                                                                                                                                                                                                      
                                ,                 	                                                                                                                        0                                                            	                                        ,                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                 	       ,                                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                                ,                                                                                                                                                                                                                            ,                                                                                             
                                                                                                                                                 ,                          	                                                                                                                                                                                                               .                                                                                                                                                                                                            #              ,                                                                                                                                                                                                                           -                                                                                                  
                                                                                                                                      ",                                                                                           *                                                                                                                                          ,                                                                                                                                                                                                                            -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                          	        ,        	                                                                                                                                                                                                                                 .                                                                                                                                                                                                            -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                           
 -                                                                                                                                                                                                                     
       ,                                                                                                                                                                                                                                      -                                                                                                                                                                                                                  
                          -                                                                                                                                                                                                                    
            -             
                                                                                                                                                                                                                
       ,                                     	                                                                                                                                                                                                     .                                                                                                                                                                                                                      	              &             -                                                                                                                                                                                                                         -                                                                                                                                                                                                                        ,               	                                                                                                                                                                                                               ,                                                                                                                                                                                                                                       	     ,                                      2                                                         
                                                                                                                                    -                                        -                                                                                                                                                                                         /                                                                                                                                                                                                                -                                                                                                                                                                                                                             ,                                                                                                                                                                                                          
                        #   
       -                                                                                                                                                                                                                                ,                                      	                                                                                                                                                                                          ,                                                                                                                                                                                                                           -                                                                                                                                                                                                                              -                   -                      
                                                                                                                                                                                                         ,                                                                                                                                                                                                                                    
       -          	      
                                                                                                                                                                                                              ,                                                                                                                                                                                                                            	       &
                   ,                                        
                                                          #                                                                                                                                         ,                                                                                                                                                                                                 	                 /                                                                                                                                                                                                                             ,                                                                                                                                                                                                             
   
                                 ,                                                                                                                                                                                                                                                 .                                                                                                                                                                                                                      .                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                          
        -           
                                                                                                                                                                                                                -                                                                                                                                                                                                                     
         -                                                                                                                                     	                                                                                         -                                                                                                                                                                                                                                        .                                                                                                                                                                                                                            
                 ,                                                                                                                                                                                                                               ,                                                                                                                                                                                                                           ,                                                                                                 	                                                                                                                                   .                                                                                                                                                                                                             
                ,                                                                                                                                                                                                                    ,                               
                                                                                                                                                                                            -                                                                                                                                                                                                                                -                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                  -                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                    	  -      	                                                                                                                                                                                                                     ,       	                                                                                                                                                                                                                                -                                      
                                                                                                                                                                                                  ,                                                                                                    .                                                                                                                                           -                                                                                                                                                                                                                                 .                                                                                                                                                                                                                                  -                                                                                                                                                                                                                                       -                                                                                                                                                                                          	                                ,                                                                                                                                                                                                                            -                                                                                         	                                                                                                                             -                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                  ,                                                                                              	                                                                                                                                              -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                 	-                                                                                                                                                                                                                                         -                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                   I                    .                                                                                                                                                                                                                                -                                                                                                                                                                                                                               -          	      	                
                                                                                                                                                                                           ,                                                                                                   	                                                                                                                                      -                                                                                               	                                                                                                                                       .                                  (                                                                                                                                                                                            -                                <                                                                                                                                                                                                  ,                                                                                                                                                                                                                     	              .                                                                                                                                                                                           	                       	         ,                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                              	             )          -                                                                                                                                                                                                                       -                                                                                                                                                                                                                              	         -                                                                                                                                        "
                                                                                              -                                                                                                                                                                                                                                 -                   ,                                     	                                                                                                                                                                                              .                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                 ,                                                                                            	                                                                                                                                -                                                                                                                                                                                                                                     .                                                                                                                                                                                                                            ,       
          	                                                                                                                                                                                                                    ,                                                                                                                                                                                                  "
                                  ,                                    
                                                                                                                                                                                              ,                                          
                                                                                                                                                                                         ,                                                                                                                                                                                                                                    %      	     ,                                                                                                                                                                                                                            #            -                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                      *        -                                                                                                                                                                                                                                          ,      	                                                                                                                                                                                                                                            ,                                                                                                                                                                                                   	                                      -                                                                                                                                                                                                                                 ,                                                                                              1                                                                                                                                            -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                             .                  -                                                                                                                                                                                                                          ,                                   	                                                   	                                                                                                                                	,                                       <                                                                                                                                                                                                       ,            	                                                                                                                                                                                                                                       ,                                        .   	                                                                                                                                                                                                   ,        
                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                    -                                                                                                                                                                                                                                  ,                                            
                                                         	                                                                                                                           
           ,                 "                                                                                                                           	                                                                                                   ,                                                                                                                                                                                                                                            ,                                                                                                                                                                                                                      ,                           	                                                                                                                                                                                                             
,         
                                                                                         -                                                                                                                                                   ,                                                                                                                                                                                                                                         ,                                     '                                                                                                                                                                                                 ,                   
                                                                                                                            	                                                                                            ,                                                                                                                                                                                                               7                                          ,                                                                                                                                                                                                                                            ,                                                                                                                                                C                                                                                                     -                                                                                                                                                                                                        & 
                          	        ,                                                                                                                                                                                                                                                    -                                                                                                                                                                                                                                        ,                
                                                                                                                                                                                                                 -                                                                                                                                                                                                                                   ,                $       	                                                                                                                                                                                                                       ,                                                                                                                                                                                                	                             ,                                                                                                                                                                                                                                  -                                                                                                                                                                                                                                -                                                                                                                                                                                                                            ,         
             	                                                                                                                  
                                                                                                     ,               
       
         
                                                                                                                                                                                                       .                                                                                                                                                                                                                                
       ,                                                                                                                                                                                                    
                                 ,                                                                                                                                                                                                                          -                                                                                                                                                                                                                                %             ,                                                                                                                                                                                                                                             .                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                            
                ,                                                                                                                                                                                                                                             -          
                                                                                                                                                                                                                              ,                                                                                                                                                                                                                          -                                                                                                                                                                                                                           	                    -                                                                                                                                                                                                                                     -                       	                                                                                                                                                                                                           ,                                                                                                                                                                                                                       ,                                                                                                                                                                                                                          "                    ,                                                                                                                                                                                                                             -                                   	   
                                                                                                                                                                                                      ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                              ,                                                                                            	                                                                                                                                      ,             .                                                                                                                                                                                                                                  .                                                                                                                                                                                                                    	              ,                                                                                                                                                                                                                            -                                                                                                                                                                                                                       !                    ,                                                                                                                                                                                                              	                                   -                                                                                                                                                                                                           
                ,          )                        	                                                                                                                                                                                                           ,                                                                                                                                           
                                                           
                                 ,                                      
                                                                                                
                                                                                                    ,                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                            ,                    
                                                                                                                             0                                                                                                  ,                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                               ,                                                                                                                                                                                                                               -               	                                                                                                                                                                                                                        ,                                  	                                                                                                                                                                                        ,             5                             	                                                                                                                                                                                                               /                                                                                                                                                                                                                                      .                                                                                                                                                                                                                                 ,                                   
                                                                                                                                                                                                 ,       	                                                                                                                                                                                                                                   ,                                                                                                                                          	                                                                                        ,                                                                                                                                                                                                                                      ,                                    
                                                                                                                                                                 !                                  ,                                                                                                                                                                                                                           ,                     	
                                                                                                                             
                                                                                                   -                                                                                                                                                                                                                             0       ,                                                                                                                                                                                                                                  /                                                                                                                                                                                                                         2               ,                                                                                                                                                                                                                                                 .                                                                                                                                                                                                                        	              #            ,                                                                                                                                           
                                                            	                            -                                                                                                                                                                                                                                           ,           	                       
                                                             	                                                                                                                                  -            
                                                                                                                                                                                                                             ,                                                                                                                                           	                                                                                         ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                     .                                                                                                                                                                                                                           #             
      ,                                                                                           
                                                                                                                               ,                                                                                                                                                                                                                                               ,        	                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                                -                                                                                                                                                                                                                         
,                    !                                                                                                                                                                                                                               -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                             -                                                                                            	                                                                                                                                        ,         
   
       *       
           
                                                                                                                                                                                                           .                                                                                                                                                                                                              #                ,                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                       -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                   ,                                 %                                                            	                                                                                                                                              ,              	       	                                                                                                                !                                                                                                     -                                      
   	                                                                                                                                                                                                  ,                                                                                                                                                                                                                                           ,                                                                                                                                                                                                          
                                   ,                 #                                                                                                                                                                                                                     ,                   %                                                                                                                                                                                                                                ,                                                                                                                                                 
                                                                                              ,                                                                                                                                        $                                                                                                     .                                                                                                                                                                                                                              ,           +                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                            -     	         
                	                                                                                                                                                                                                        ,                
                                                                                                                                                                                                                ,                   0       
                                                                                                                                                                                                                ,                                                                                               	                                                                                                                               	     
    ,        
                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                  -                                                                                                                                
                                                                                          ,                                                                                                                                                                                                                      /                                                                                                                                                                                                                      	      ,                                                                                                                                                                                                                          	                -                                                                                                                                                                                                                                     ,                                                                                                	                                                                                                                                 .                                                                                                                                                                                                                                 	      ,                                                                                               	                                       
                                                                                         -                                	                                                                                                                                                                                                    ,                                 	                                                                                                                                                                           	              -                                                                                                                                                                                                                                   ,                                                                                                                                        	                                                                                     ,                                                                                                                                                                                                                          ,                                                                                                                                                                                                                 .                                                                                                                                                                                                            	      	           .                                                                                                                                                                                                                         -                       	                                                                                                                                                                                                                -                                                                                                                                                                                                                                  
    ,                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                           /           
    ,                    3                                                                                                                                                                                                                         -             
                                                                                                                                                                                                            ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                  B                ,                                                                                                                                         
                                                                                               -             
                                                                                                                                                                                                            ,                                                                                                                                                                                                                                       ,                                                                                                                                                                                                               
                          
,                                                                                                      	                                                                                                                             2           	     .                                                                                                                                                                                                                           -                                    /                                                                                                                                                                                                        ,                                                                                                                                                                                                                                               ,                                                                                                                                                  
                                                                                             .                                                                                                                                                                                                                                   /                                                                                                                                     )                                                                                                    ,                                                                                                                                                                                                                                  ,          -                                                                                                                                                                                                                                   .                                                                                                                                                                                                                           ,                                                                                                                                      	                                                                                          .                                                                                                                                                                                                                              !            .                                       	                                                                                                                                                                                      	             -                                                                                                                                                                                                                            -                                                                                                                                                                                                                               .               	     	                                                                       	                                                                                                                               	            -                                                                                                                                                                                                                                    .                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                 ,                	                                                                                                                                                                                                                       ,                   
                                                                                                                                                                                                              ,                                                                                                                                                                                                                                  
        .                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                          -              	                                                                                                                                                                                                                  -                                                                                                                                                                                                                
                -                                                                                                                                                                                                                              
   ,                                                                                                                                                                                                                               #          
     ,        
                                                                                                                                                                                                                            -                                                                                                                                                                                                                       -                                                                                                                                                                                                              	               .                                                                                                                                                                                                                               ,       	                	             	                                                                                                                                                                                              -                                                                                                                                                                                                                -              	                                                                                                                                                                                                      
     ,                                         
                                                                                                                                                                                                     ,                      
                                                                                                                                                                                                        .                                                                                                                                                                                                                         
      "       ,             %       
                                                                                                                                                                                                               ,                                                                                                                                                                                                                                      -              &                                                                                                                                                                                                 	                   .                                                                                                                                                                                                                                         -                                                                                                                                                                                                                                   -                                                                                                                                                                                                                                       -                                                                                                                                                                                                                                           .                                                                                                                                                                                                                         ,                                                                                           
                                                                                                                             ,                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                              
         	      -                                                                                                                                                                                                                                    -                                                                                                                                                                                                                                          ,                    !                                                                                                                                                                                                                     ,                                                                                                                                                                                                      	                              	   -                                                                                                                                                                                                                         -                                                                                                                                     	                                                           
                                     ,                         
                                                                                                                                                                                                              -                                                                                                                                                                                                                                   .                                                                                                                                                                                                                                 	    .                                                                                                                                                                                                                        ,                 '                                                                                                                       
                                                                                                  ,          	             
                                                                                                                                                                                             
                 -                  
                                                                                                                                                                                                         0                  -                                                                                                                                                                                                                        -                                                                                                                                   
                                                                                                 .                                                                                                                                                                                                                                   .                                                                                         
                                                                                                                                 ,                                  	                                                                                                                                                                                                  ,                                                                                                                                                                                                  '                                   .                                      
                                                                                                                                                       	                                  ,                                                                                                                                                                                                                      .                                                                                                                                                                                              	                                   ,                                                                                                                                                                                                       	  	                             .                                                                                                                                                                                                                         ,                                                                                                                                                                                                                         .                                                                                                                                                                                                                                    
      -                                                                                                                                                                                                                         -               	                                                                                                                                                                                                         	             .                                                                                                                                                                                                                         	-                                                                                                                                                                                                                           
                    -                                                                                                                                                                                                                           ,                       
          	                                                                                                                                                                                               ,                                                                                                  
                                                                                                                                -                                                                                                                                                                                                                     "	              ,                                                                                                                                                                                                                               /                                                                                                                                                                                                                      ,                                                                                                                                                                                                                         -                                                                                                                                                                                                                              .               	         	                                                                                                                                                                                            .                                                                                                                                                                                                                                -                                                                                                                                                                                                                           ,                	                                                                                                                                                                                                                  ,                                                                                           
                                                                                                                                .                                                                                                                                                                                                                                   -                                                                                                                                                                                                                                -     	                                                                                                                                                                                                                              ,                                                                                                                                                                                                                         -                                                                                            	                                                                                                                                     .                                                                                                                             	                                                                                      .                                                                                                                                                                                                                                    ,                                                                                                                                                                                            	                                 	,                                                                                                                                                                                                   
                                 .                                                                                                                                                                                                                        .                                                                                                                                                                                                	                                         .                                                                                                                                                                                                                           .         .       %                                                                                                                                                                                                                        -                                                                                                                                                                                                                          	      -                                                                                                                                                                                                                                   ,                                                                                   	                                                                                                                             	    -                                                                                                                                                                                                                                 /                                                                                                                                                                                                                 	       .                                                                                                                                                                                                                              ,               
                                                                                                                                                                                                                       ,                	                                                                                                                                                                                                      ,                                                                                                                                                                                                                        -                
                  
   
                                                                                                                                                                                                   .                                     	                                                                                                                                                             %                            .                                                                                                                                                                                               	                                     -                                                                                                                                                                                                                    .                                                                                                                                                                                                                              '       
      ,                                                                                                                                                                                                                              )                .      	 	               	                                                                                                                                                                                                                   ,                                       	   
                                                                                                                                                                        
            .                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                 -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                          
           /                                                                                                                                                                                                                                       
     -                                                                                                                                                                                                                                ,                                  
                                                                                                                                                                                              /                                                                                                                                                                                                                       -                                                                                                                                                                                                                     $           	      -                                                                                                                                                                                                                           	,                                                                                                                                                                                                                                     -                                                                                                                                                                                                                   ,                                                                                                                                                                            
                                                           ,                                                                                                                                                                                                                                /                                                                                                                                                                                                                                 	             -                                                                                                                                                                                                                        .                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                              -        	                 
                                                                                                                                                                                                                   ,                                                                                                                                                                                                                            -                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                   ,                                 	                                                                                                                                                                                                    -                                                                                                                              	                                                                                       /                                                                                                                                                                                                                         ,                                                                                              	                                                                                                 	                     
        ,                                                                                                	                                                                                                                                    -                             	                                                                                                                                                      	                                    -                                                                                                                                                                                                                     
-                                                                                                                                                                                                                                        .                                                                                                                                                                                                                          	            -                                                                                                                                                                                                 	                                ,                                                                                                                                                                                                                                      -                                                                                                                                                                                                                 	                 -                                                                                                                                                                                                                                        /                                                                                                                                                                                                                            ,                                                                                                                                                                                                                     	                    /                                                                                                                                                                                                                   .                                                                                          
                                                                                                                                            ,                                                                                                                                                                                                                     ,                                                                                                                                                                                                                    -                                                                                                                                                                                                                           ,                                                                                                                                                                                                                        ,                                                                                                                                                                                                                          -                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                      .                                                                                                                                                                                                                        ,               
                                                                                                                                                                                                             -                                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                        .                                                                                                                                                                                                                    .           
                                                                                                                                                                                                      
                         -                                                                                                                                                                                                                   -                                                                                                                                                                                                                    
               /                                                                                                                                                                                                               	.                                                                                                                                                                                                                                                 ,                                                                                                                                                                                                  
                              /                                                                                                                                                                                                                 .                                                                                                                                                                                                                           ,                          
                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                  4                   ,                                                                                                                                                                                                                                       -                                                                                                                                                                                                                         -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                              0             	       .           
                                                                                                                                                                                                                      	/                                                                                                                                                                                                                           ,             	                                                                                                                                                                                                          ,                                                                                                      
                                                                                                                                        -                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                           .                                   *                                                                                                                                                                                             ,                                                                                                                                                                                                                                       
      ,                                                                                                                                                                                                                               -                                                                                                                                                                                                                               -                                                                                                                                           -                                                                                                 ,                                                                                                                                                                                                            	                           .           .                     
                                                                                                                                                                                                          -                                                                                                                                                                                                                                -              	                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                          3             .                     
                                                                                                                                                                                                                .                                                                                                                                                                                                                
    ,          )                                                                                                                                                                                                                 	                 -                                                                                                                                                                                                                             ,                                                                                                                                
                                                                                          -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                        
  .                                                                                                                                                                                                                                           -                                     
                                                                                                                                                                                             ,                                                                                                                                                                                                                              
-                                                                                                                                                                                                                                        ,                                                                                                	                                                                                                                                  -                                                                                                                                                                                                                    	                     ,                                                                                                                                             
                                                                                             ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                9                                       -                                                                                                                                                                                                                               0      
       ,                                                                                                                                                                                                                                      .                     
                                                                                                                                                                                                        $      
      -                                                                                                                                                                                                                           ,        
                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                     !                  ,                                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                           -                                                                                                                                                                                                                         -                                                                                                                                                                                                                      
     ,                                                                                                                                                                                                                                           N             ,                                                                                                                                      	                                                                                                 -                                                                                                                                                                                                                                 <            ,            	                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                           	      ,               (                                                                                                                                                                                        
                                        ,                                                                                                
                                                                                                                                     ,                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                "             "      ,                                                                                                  +                                                                                                                                                     ,                                       =                                                                                                                                                                                                       -                                
                                                                                                                                                                                ,                                                                                                                                                                                                              	                              ,                                                                                                                                                                                                            4                                     	,                                                                                                                                                  0                                                           
                                 ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                             .             ,            
      	                                                                                                                                                                                                                            -                                                                                                                                                                                        
                                 -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                         =             ,            (                                                                                                                                                                                                                                 .                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                 -                                                                                                                                                                                                                              	      +             ,                                                                                                                                                                                                                                                ,                                                                                          	                                                                                                                                      ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                  
                                 ,                      
         
                                                                                                                                                                                                    ,                                                                                                                                                                                                                     	      .                                                                                                                                                                                                                          )            ,                                                                                                                                                                                                                        
                -          
                                                                                                                         
                                                                                              ,                                      
                                                                                                  	                                                                                    .                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                #        ,                                                                                                                                                                                                                                   +             -                                                                                            	                                                                                                                                        .                                                                                                                                                                                                                                  5      	      .                                                                                                                                                                                                                               -                                                                                                                                                                                                                                   ,                                                                                                                                  
                                                                                             -                                                                                                                                                                                                                            6             ,                                     1                                                                                                                                                                                               -                                 +                                                          	                                                                                                                                       /                                                                                                                                                                                                                       /
                                                                                                                                                                                                                                 -                                                                                                                                                                                                                            /                                                                                                                                                                                                             ,                                                                                                   	                                                                                                                               -                                                                                                                                    	                                                                                              0             #                                                                                                                                                                                                               ,                                                                                                                                            	                                                                                         /                                                                                                                                                                                                                        /            
                                                                                                                                                                                                                    /                                                                                                                                                                                                                          ,                                                                                                                                      	                                                                                             0                                                                                                                                                                                                                       ,                                      
                                                                                                                                                                                                ,                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                              -                                                                                                                                                                                                                                      /                 
                                                                                                                   
                                                                                                ,                                                                                                                                                                                                                                            ,                 	                                                                                                                                                                                        "                              
          0                                                                                                                                                                                                                           -                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                       
        ,                                                                                                                                                                                                                                                   /                                                                                                                                                                                                                              ,                                                                                                                                                                                                                          -                                                                                                                                        
                                                                                      -              	      
                                                                                                                                                                                                     .                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                 /                                                                                                                                                                                                                  -                                                                                                                                                                                                           /                                                                                                                                                                                                                   	 /                                                                                                                                  	                                                                                       .                                                                                                                                                                                                                 0               
                                                                                                                                                                                                   0                                                                                                                                                                                                        	      1                                                                                                                                                                                                           .                                                                                                                                                                                                             .      	                                                                                                                                                                                                       1                                                                                                                                                                                                             2                                                                                                                                                                                                                        0                                                                                                                                                                                                                        .                                                                                                                                                                                                                  3                                                                                                                                                                                                              1       	                                                                                                                                                                                                     .                                                                                                                                                                                                                  /                                                                                                                                                                                                                     /                                                                                                                                                                                     
                        ,    	         	                                                                                                                                                                                                             .           
                                                                                                                                                                                                                     -                                                                                                                                                                                                                   ,                                                                                                                                                                                                                 /     
    	                                                                                                                                                                                                                     ,                                                                                                                                                                                                                            "	             -                                                                                                                                                                                                                           -                                                                                           
                                                                                                                                .                                                                                                                                                                                                            -                                                                                                                                                                                                                -                                                                                                                                                                                                                          .                                  

                                                                                                                                                                                        /                                                                                             	                                                                                                                             -                                                                                                                                                                                                              /                                                                                                                                                                                                         /                                                                                                                                	                                                                                  /                                                                                                                                                                                                                  .                                                                                                                                                                                              	                             ,                             	                                                                                                                                                                                              /                                                                                                                                                                                                                  .                                                                                                                                                                                                              0                                                                                                                                                                                                                       
                  /                                                                                                                                                                                                             -                                                                                                                                                                                                                  -               
                                                                                                                                                                                                                 1                                                                                             	                                                                                                                             .                                                                                                                                                                                                                       .                                                                                              
                                                                                                                          -   	                                                                                                                                                                                                                               /                                                                                                                                                                                      	                             
    /            	                                                                                                                                                                                                    /                                                                                                                                                                                                               
     /           	                                                                                                           
                                                                                         ,                              	                                                                                                                                                                                            .                	                                                                                                                                                                                                           .                                                                                                                                                                                                                    1                                                                                                                                                                                                                     	    /                                                                                                                                                                                                               -         
                                                                                                                                                                                                      	          -                                                                                                                                                                                                                   .                                                                                                                                                                                                                                        /                                                                                                                                                                                                                       0                                                                                                                                                                                                                  .                                                                                                                                                                                                       -                                                                                                                                                                                                                /                                                                                                                                                                                                             .                                	                                                                                                                                                                                          0                                                                                                                                                                                                      ,       
      	                                                                                                                                                                                                               .                                                                                                                                                                                                                                  .                                                                                      
                                                                                                                              /                                                                                                                                                                                                                ,   	                                                                                                                                                                                                                          ,                                                                                                                                                                                                                           )	               ,                "                                                                                                                       
                                                                                             .                                                                                                                                                                                                                            .     
                                                                                                                                                                                                              0                                                                                                                                                                                                         -                                                                                                                                                                                                                              /                                                                                                                                                                                                                      1                                                                                                                                                                                                                 2                                                                                                                                                                                               	0                                                                                                                                                                                                            1                                                                                                                                                                                                                   1                                                                                                                                                                                                         .                                                                                                                                                                                                                             ,           "                      
                                                                                                                                                                                                     -                                                                                                                                                                                                                    .        
   
                                                                                                                                                                                                            .                                                                                                                                                                                                                
       	                /           	                                                                                                                                                                                                          /                                                                                                                                                                                                                   .                                                                                                                                                                                                                                 /             	                                                                                                                                                                                                            ,                                                                                                                                                                                                                      /                                                                                                                                                                                                                             /                   	                                                                                                                                                                                                          /                                                                                                                                                                                              	                          	   .                 	                                                                                                                                                                                                         -                                                                                                                                                                                                                
                 	  -              
                                                                                                                    
                                                                                        .                                                                                      
	                                                                                                                               0                                                                                                                                                                                                            	                  ,                                                                                                                                                                                                                             5                                                                                                                                                                                                                1                                                                                                                                                                                                         /                                                                                                                                                                                                                        .                                                                                                                                                                                                            
               	  3                                                                                                                                                                                                                   /                                                                                                                                                                                                                        -                                                                                                                                                                                                                          -                                                                                                                                                                                                             	       /                                                                                                                                                                                                                /                                                                                                                                                                                                                 -                                   	                                                    
                                                                                                                                       1                                                                                                                                                                                
                       -                                                                                                                                                                                                                        .                                                                                                                                                                                                                                -                                                                                                                                                                                                                .                                                                                                                                                                                                                  -         	                                                                                                                                                                                                              .                                                                                                                                                                                                                       $            -                                                                                                                                                                                                                       /                                                                                           	
                                                                                                                                 .                          
                                                                                                                                                                                        .                                                                                     	                                                                                                                              ,                                 
                                                                                                                                                                                              -                              
                                                                                                                                                                                      /                                                                                                	                                                                                                                           .                                                                                                                                                                                                     1                                                                                                                                                                                                                 /                                                                                                                                                                                                                  .                                                                                                                                                                                                           .                                                                                                                                                                                                                         
   -                                  	                                                                                                                                                                                               /                                                                                                                                                                                                                     /                                                                                                                                                                                                                .                                                                                                                                                                                                           
                        0                                                                                                                                                                                                                   -                                                                                                                                                                                                                    ,   	   	                                                                                                                                                                                                                            /                                                                                                                                                                                                                            ,                                                                                                                                                                                                                 .                                                                                                                                                                                                                  	                ,   	               	                                                                                                                                                                                                                  -                                                                                                                                                                                                      	                         ,                                                                                                                                                                                     
                              ,                                                                                                                                                                                                                                	.                                                                                                                                   
                                                                                           .                                                                                                                                                                                                                                	 ,                                                                                                                                                                                                                     	       -                                                                                                                                                                                                                    
-                                                                                                                                                                                                                      ,                                                                                                                                                                                                             ,                                                                                                                                                                                                                                            -        #                                                                                                                                                                                                                 /                                                                                                                                                                                                                               ,                                                                                               
                                                                                                                                -                                    
                                                                                                                                                                              	           -                                                                                                                                                                                                                       ,                                                                                                                                                                                                              
               ,                                 	                                                                                                                                                            	                                    .                                                                                                                                 	                                                                                            ,                                                                                                                                                                                                                                      
-                                                                                                                                   
                                                                                             ,            	                                                                                                                                                                                              	                  .                     
                                                                                                                                                                                                  	           -                                                                                                                                                                                                                     -                                                                                                                                           
                                                                                    	,                                                                                                                                                                                                                                       ,          	                                                                               	                                                                                                                                   .                                                                                       
                                                                                                                             ,           	                                                                                                                                                                                                               ,                                                                                               
                                                                                                                                    ,                                                                                          
                                                                                                                                
-                                                                                                                                                                                                                                     ,                                 	                                                                                                                                                                                        -                                                                                                                                                                                                                                .                                                                                                                                                                                                                           
,                 
                                                                                                                                                                                                               ,                                                                                                                                                                                                                        ,                                                                                                                                                                                                                    ,           	                                                                                                                                                                                                             -                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                        
       .                     
                                                                                                                                                                                                     .                                                                                                                                                                                                  	             ,                                                                                                                                                                                                                                   -                                                                                                                                                                                                                           ,           
                                                                                                                                                                                                              ,     
                         	                                                                                                                                                                                   
               ,                                                                                                                                                                                                                                     	-                                                                                                                                                                                                                                        .                                                                                                                                                                                                                               ,                                                                                                                                                                                                      	                             -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                         	-                                                                                                                                                                                                                                  -                               	                                                                                                                                                                                           .                   
                                                                                                                                                                                                                       	     ,                                                                                                                                            	                                                       	 	               
                -                                                                                                                                                                                                                                            -                               
                                                                                                                                                                                               -                                                                                                                                                                                                                                        .                                                                                                                                                                                                                              -                                                                                                                                                                                                                              -                                                                                                                                                                                                         		               -                                                                                                                                                                                                                          (                 ,                                                                                                                                                                                                                                 0                                                                                                                                                                                                                 ,                                                                                                                                                                                                         
                            .                	       	                                                                                                                                                                                                                -                                                                                                                                            
                                                                                           ,                  %                                                                                                                                                                                                                        .                                                                                                                                                                                                                       
     ,                                                                                                                                    
                                                                                  ,                                                                                                                                                                                                                     
             
        ,                                                                                                                                       
                                                                                              -                                                                                                                                                                                                                              	      -                                                                                                                                                                                                                             -                                                                                                                                                                                                                                        -                                                                                                
                                                                                                                                ,                                                                                                                                                                                                                                         -                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                            
         
     ,                                                                                                                                                                                                    	                            
    ,                                                                                                                                                                                                                                              -                                   	                                                                                                                                                                                                     ,                                                                                                                                                                                                                                          $            .        	                                                                                                                                                                                                                            ,                                      
                                                                                                                                                                                   -                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                   ,            '              
                                                                                                                                                                                                                    .                                                                                                                                                                                                                               ,      	                                                                                                                                                                                                                      -                                                                                                                                                                                                                             ,         	                                                                                                                                                                                                                          -                                                                                                                                                                                                                                "     
       ,       	  !                                                                                                                                                                                                                       -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                   .                                                                                                                                                                                                                             -                                                                                                                                                                                                                 .                                                                                                                                                                                                                                   ,              	                                                                                                                                                                                                        ,             	                                                                                                                                                                                                      .                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                    /                                                                                                                                                                                                                            .                                                                                                                                                                                                                                     -                                                                                                                                                                                                                              -                                                                                                                                                                                                               	-            	    
                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                  	     
/                                                                                                                             
                                                                                              ,                                                                                                                                                                                                
                        	-                                                                                                                                                                                          
                                    .                                                                                                                                                                                                             
                        ,                                                                                                                                                                                                                                               -                                                                                                                                                                                                                	  -                                                                                                                                                                                                             .                                     	                                                          
                                                                                                                                           ,                 
                     	                                                                                                 
                                                                                             /                                                                                                                                                                                                                       ,                         	                                                                                                                                                                                           ,                                                                                                    	                                                                                                   
                 	        -                                                                                                  
                                                                                                                                  .             
                                                                                    	                                                                                                                                           ,                                                                                                                                                                                                                             ,                                                                                                                                                                                         	                          ,                                                                                                                                                                                                                                     
.                                                                                                                                                                                                                                        -                                                                                                                                                                                         
                                  ,                                                                                                                                                                                                                                  &         -                
                                                                                                                     	                                                                                            .                                                                                                                                                                                                
                                -                                                                                                                                                                                                                   -                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                          -                                                                                                                                                                                                                   )              .       	                                                                                                                                                                                                                 ,                                                                                                     
                                           	                                                                          	              -                     	                                                                                                                                                                                                              ,                                                                                                                                                                                                                                 
   ,        
      
                
   	                                                                                                                                                                                              ,                                                                                                                                                                                                                               ,                                                                                                                                                                                                             
           .                                                                                                                                                                                                                      -                                                                                                                                                                                                                                      -                                                                                                                                                                                                                         ,                                                                                                                                                                                                                 
            -                                                                                                                                                                                                                              0                       	                                                                                                                                                                                                    ,                                                                                                   	                                                                                                                           .                                                                                                                                                                                                                                         ,                                                   	                                                                                                                                                                      -                      
                                                                                                                                                                                                     
   ,                                                                                                                                                                                                          
                  ,         	             	           	                                                                                                                                                                           
                  -                                                                                                                                                                                                                            -                  
                                                                                                                                                                                                     	      .                                                                                                                                                                                                                    .                                                                                                                                                                                                            -                                                                                                                                                                                                               	            ,                                                                                                                                                                                                                                          -                                                                                                                                                                                                           	                /          	                                                                                                                                                                                                                 1                                                                                                                                                                                                                  	   ,                                                                                                                                                                                                                                ,                                                                                                                                                                                                                               /                                                                                                                                                                                                                    -                                                                                              
                                                                                                                            .                                                                                                                                                                                                                           	/                                                                                                                                                                                                                 .                                                                                                                                                                                                               -                                                                                                                                                                                                              .                                                                                                                                                                                         
                                   ,                                                                                                                                                                                                  
                        ,                                                                                                                                                                                                                                            0                                                                                                                                                                                                       .                                                                                                                                                                                                                            .                                                                                                                                                                                                                                  ,                                                                                                                                                                                                 	                                .                                                                                                                                                                                                                        ,                                                                                                                                                                                                                           -                                                                                                                                                                                                   	                       #   	     0                                                                                                                                                                                                                             .                                                                                                                                                                                                                          -                                                                                                                                                                                                                            1                                                                                                                                                                                                                      ,          	                       	                                                                                                                                                                                              ,                                                                                                                                                                                                                                    -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                             '                                 .                                                                                                                                                                                                                                	           .                                                                                                                                                                                                                        
      -                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                            -                                                                                                                                                                                                               
     
        ,           
       
                     	                                                                                                  	                                                                                                -                 	                                                                                                                                                                                                                  .                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                      (   	      ,                                                                                          
                                                                                                                              -            
                                                                                                                                                                                                                        -                                                                                                   	
                                                                                                                                
     ,                        
         
                                                                                                                                                                                                 ,                                                                                                                                                                                                                           
     .                                                                                                                                                                                                                                !           -                                       +                                                                                                                                                                                                            ,                                      4                                                                                                                                                                                                             -                                	                                                                                                                                                               	                                  ,           !                                                                                                                                                                                                                                   .                                                                                                                                                                                                                        ,                         
                                                                                                                                                                                                       .                                                                                                                                                                                           
                              ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                       $             ,                6                                                                                                                         	                                                                                                  ,                                                                                                                                                                                                                                 -                               	                                                                                                                                                                                            ,                                                                                                                                                                                                                                       ,       
                                                                                      "                                                                                                                                                  ,                                                                                                                                                                                                                                                 ,                                  )                                                                                                                                                                                                         ,                                                                                                                                                                                                                               ,                                                                                                                                                
                                                                                    	      -                         	                                                                                                                                                                                
                                        ,                                                                                                                                           1                                                                                                    ,                                                                                                                                                                                                                                   #   	       -               	                                                                                                                                                                                                                               .                                                                                                                                                                                                                   
           	    -                                                                                                                                                                                                                       -                                                                                                                                                                                                                             ,            &                         	                                                                                                                                                                                                           .                                                                                                                                                                                        	                             ,                                                                                                                                                                                                                 
                .                                                                                                                                                                                                                                  ,                                                                                                                                           
                                                           	                          	       /                                                                                          	                                                                                                                                           ,                               *                                                                                                                                                                                                   .                                                                                                                                                                                                                                )        ,                                                                                                                                                                                                                              -                               	                                                                                                                                                                                     .                                                                                                                                                                                                                         	,                                                                                        	                                                                                                                           ,                                                                                                                                                                                                                                          ,           	                                                                                                                            	                                                                                        .           	                                                                                                                                                                                                                   
  ,                                                                                                                                     	                                                                                     -                                                                                                                                                                                                                        
              ,                                    
   
                                                                                                                                                                               	            .     
                                                                                                                                                                                                                   -                                                                                              
                                        	                                                                                            ,                                                                                                                                  		                                                                                           /                                                                                                                                                                                                        -         
                                                                                                                                                                                                                 ,                                    
                                                                                                                                                                                   	          .                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                            ,                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                     ,          	     	                                                                                                                                                                                                                           /                                                                                                                                                                                                                         ,                                                                                                                                    
                                                                                         ,                                                                                                                                                                                                                                  $          
 ,   	                                                                                                                                                                                                                                   /                                                                                         	                                                                                                                                   ,                                                                                                                                                                                                                          -                                                                                                                                                                                                                    
     -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                         -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                                 -                                                                                           	                                                                                                 
                                     ,                                                                                                                                                                                                                                          ,                                                                                                                                          
                                                         
                                      ,                                                                                                                                                                                                                       ,               		                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                                -          !                                                                                                                                                                                                                          /                                                                                                                                                                                                                       -                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                 -                                                                                                                                                                                                                                         /                                                                                                                                                                                                                         -                                                                                                                                                                                                                                -                                                                                                                                                                                                       
                             
        ,                                                                                                                                    
                                                                                              -                                                                                                                                                                                            
                               ,                                                                                       
                                                                                                                                  -                                                                                                                                                                                                                                             -                                                                                                                                                                                                                                    -                                                                                                                                  	                                                                                      -                                                                                                                                                                                                                          
    -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                       	      
               ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                                           -                                                                                                                                                                                                                         	     ,                                                                                                                                                                                                                     .                       	                                                                                                                                                                                               	       ,                                                                                                                                                                                                                                        ,           (                                                                                                                                                                                                                       ,                                                                                                                                                                                                            (                                  ,                                                                                                                                                                                                                                          ,             	                                                                                                                                                                                                               ,                                                                                                                                              	                                                                                      .                                                                                                                                                                                                                     -                                                                                                                                     	                                                                                        ,                                                                                                                                                                                                                                     -                                                                                                                                      	                                                                                     /                                                                                                                                                                                                                 .                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                 -                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                             -       	                                                                                    	                                                                                                                                           ,                                                                                                                                                                                                                                 	,                                                                                                                                                                                                                                      ,                                                                                                                                           #                                                                                                   ,                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                   
       -     	                                                                                                                                                                                                                            .                                                                                                                                                                                             
 	                           ,                                                                                                                                                                                                                                        -                                                                                                                                                                                                                        #        -          $                                                                                                                                                                                                                               .                             
                                                                                                                                                                             0               	                                                                                                                                                                                                               1                                                                                                                                                                                                                    ,                  
       
                                                                                                                                                                                                         .                                                                                  
                                                                                                                                    ,                                   (                                                                                                                                                                                                 ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                    -                                                                                                                                                                                                                            ,                                                                                                                                                                                                                         -                                                                                                                                                                                                                                    -                                                                                                                                                                                                           .                                                                                                                                                                                                                          	       
   /                                                                                                                                                                                                                  -                                                                                                                                                                                                                                        .                                                                                                                                                                                                                  .                                                                                                                                                                                                                	             ,                                                                                                                                                                                                                                 .                                                                                                                                                                                                                             -                                                                                                                                                                                                                  	.                                                                                                                                                                                                                              ,                                                                                                                                                                                                  	                               ,                                                                                                                                                                                                                             -                                                                                                                                                                                                 	   
                          
        ,                                                                                                                                            *                                                                                                 ,                                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                     .                                                                                                                                
                                                                                            ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                   -                ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                       .                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                          ,                                         	                                                        2                                                                                                                                                 ,                                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                	           ,                                                                                                                                         '                                                                                                -                 
                                                                          
                                                                                                                                  ,                                                                                                                                                                                                                                         (        ,                                                                                                                                                                                                    
 
                                   -                                                                                                                                                                                                                        -                                                                                                                                                                                                                              .                                                                                                                                                                                                                                     ,           $           
                                                                                                                                                                                                           -                                                                                                                                                                                                               -                                                                                                                                                                                                                   ,                                                                                                      
                                                                                                      	                             ,                                    
                                                                                                                                                                                  /                                                                                                                                                                                                                       ,                                      
                                                                                                                                                                                                    ,                                                                                                                                                                                              
                                   ,                                                                                                                                                                                                                            .                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                      -                       
                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                          	        	   ,                                                                                                                                                                                                                           -                                                                                                                                                                                                                                         .                                                                                                                                                                                                                  -                                                                                                                                                                                                                       
                 ,                                                                                                                                                                                                                 	             -                                                                                                                                                                                                                  
                 ,                                                                                        	                                                                                                                    .            
                                                                                                                                                                                                                 	          ,                                                                                                                                                                                             
                          	   .                                                                                                                                
                                                            	                                     ,                                                                                                                                                                                                                                       ,                                                                                                                                                                                                         	                                  ,                                                                                                                                                                                                                        		     !          ,                   &                                                                                                                                                                                                                                  .                                                                                                                                                                                                                            .                                                                                                                                    	                                                                                        ,                                     
                                                         
                                                                                                                           )                  ,                 *                                                                                                                      	                                                                                                      /                                                                                                                                                                                                                          -                           	                                                                                                                                                                                               ,                                                                                                

                                                                                                                                    -                                                                                                                                                                                                                   	                ,                                                                                                                                                                                                                                          ,          
                                                                                                                                                                                                                         ,                                                                                                                                                                                                                             
      ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                   
     ,                         	              
                                                                                                                                                                                              ,                                                                                                                                                                                                                       
,              	                                                                                                                       !                                                                                                   .                                                                                                                                                                                                                              ,             #       	                                                                                                                                                                                                                                  0                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                   .                                                                                         
                                                                                                                   
              ,                   	                                                                                                                                                                                                               ,                                                                                                                                                                                                                                   -         
                                                                                                                                                                                                                         -                                                                                                                                                                                                                             ,                                                                                                                                                                                                                          ,                                                                                                                                                                                              
                           ,                                                                                                                                                                                                                            ,                                                                                        	                                                                                                                                        -          
                                                                                                                                                                                                                       .                     	                                                                                                                   
                                                                                      /         	                                                                                                                                                                                                                   ,                                                                                              
                                                                                                                                -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                                   	    -                                                                                             
                                                                                                                 	                   -                             	                                                                                                                                                                                                 .                                                                                                                                                                                                                     ,                                                                                                                                                                                                                           
          ,                                                                                                                                                                                                            
              ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                        
   -          
   	                                                                                                                                                                                                        ,                                                                                                                                                                                                                               
    ,                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                          
           -             
                                                                                                                                                                                                         	          ,                                                                                                                                                                                                                                 #               ,                        
                                                                                                                                                                                                          .                                                                                                                                                                                                                
             -       	   
                                                                                                                                                                               	                                ,                                                                                                       	                                                                                                                                    
  ,                                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                        
               .            	                                                                                                                                                                                                                     ,                                                                                                                                                                                                          
                              ,                                                                                                                                                %                                                                                                ,                                                                                                                                         
                                                                                   	          ,                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                      4   	   
     -                                                                                                                                                                                                                                       .                                                                                                                                                                                                                        -                                                                                                                                                                                                                         ,                                                                                                                                                                                                                            
     ,                                                                                                                                                                                                                                         -                                                                                                                                                                                                                
     -                                                                                                                                                                                                                            ,                                                                                                                                                                                                                   !   	         ,          
                                                                                                                                                                                                                            ,           	                                                                                                                                                                                                                       
      ,                                                                                                                                                                                                                           	          /                                                                                                                                                                                                             -                                                                                                                                                                                                                             -                                                                                                                                                                                                                   1                                                                                                                                                                                                                         ,                                                                                            
                                                                                                                                       -    	 	                           	                                                                                                                                                                                                      -                                                                                                                                                                                                                                 /                                                                                                                                                                                                                                  -                                                                                                                                                                                                               
           .                                                                                                                                                                                                                         0                                                                                                                                                                                                                  	 -                                                                                                                                                                                                                        	         /                                                                                                                                                                                                                -                                 	                                                                                                                                                                                          ,                                                                                                                                                                                                          !             1                                                                                                                                                                                                                             0                                                                                                                                                                                                                      /                                                                                                                                                                                                                      /                                                                                                                                                                                                                    .                                                                                                                                                                                                                  -                                                                                                                                                                                                                                   -                                                                                                                                                                                                             .                                                                                                                                                                                                              .   	                                                                                                                                                                                                                          .                                                                                                                                                                                                                   #                ,                                                                                      
                                                                                                                          ,                                                                                                                                                                                                              ,   	  	                                                                                                                                                                                                                    /                                                                                       
                                                                                                                            	.  	                                                                                                                                                                                                              -                                                                                                                                                                                                                    /                                                                                                                                                                                                                   /                                                                                                                                                                                                     -                                                                                                                  
                                                                                        /                                                                                                                                                                                                        .                                                                                                                                                                                                                        -                                                                                                                                                                                                                              ,          	                                                                                                                                                                                                             .                                                                                                                                                                                                                              /           	                                                                                                                                                                                                             -           
                                                                                                                                                                                                                      0                                                                                                                                                                                                                .                                
                                                                                                                                                                               /     	                         	                                                                                                                                                                                     -                                                                                                                                                                                                                      /                                                                                                                                                                                                                   .                                                                                         	                                                                                                                                  .                                                                                                                                                                                                                          /                                                                                                                                                                                                          
       .                                                                                                                                                                                          	                              ,                                                                                                                                                                                                                	        .                                                                                                                                                                                                                       -          	                              	                                                                                                                                                                                             .         	                                                                                                                                                                                                                      ,                                                                                                                                                                                                              
                -                       	                                                                                                                                                                                                             ,             	                                                                                                                                                                                                   
       -                                                                                                                                                                                                                 -                                                                                                                                                                                                                   ,                                                                                                                                                                                                                          /                                                                                                                                                                                                              -                                                                                                                                                                                                                       .                                                                                                                                                                                                                %          .                                                                                                                                                                                                                                /                                                                                                                                                                                                                       ,                                                                                                                                                                                                                         .                                                                                                                                
                                                                                         -         	            	                                                                                                                                                                                             /                                                                                                                                                                                                                              .                                                                                                                                                                                                                     -                                                                                                                                                                                                       
          /                                                                                                                                                                                                                      /                                                                                                                                                                                                                %                 -                                                                                                                                                                                                                     /                                                                                                                                                                                                                .    	                                                                                                                                                                                                            0                                                                                                                                                                                                                     .                                                                                                                                                                                                                              .                                                                                                                                                                                                  
              .                                                                                                                                                                                                                          .                                                                                                                                                                                                          -                                                                                                                                                                                                            /                                                                                                                                                                                                              0                                                                                             	                                                                                                                    .                                                                                                                                                                                                          
                    -                                                                                                                                                                                     
                             .                                                                                                                                                                                                           	           .          
                                                                                                                                                                                                           .         	                                                                                                                                                                                                                    .                                                                                                                                                                                                                   0                                                                                                                                                                                                                  .                                                                                                                                                                                                                   1                                                                                                                                                                                                                  ,                 	                                                                                                                    
                                                                                      .                                                                                                                                                                                                                               .                                                                                                                                                                                                            /                                                                                                                                                                                                              	 
       -                                                                                                                                                                                             
                              .                                                                                                                                                                                                                   .              	                                                                                                                 	                                                                                            -                                                                                                                                                                                                                            .                                                                                                                                                                                                                            ,                                                                                                                                                                                                                            .                      	                                                                                                                                                                                                            ,                                                                                                                                                                                                                      -                                                                                                                                                                                                                       /                                                                                                                                                                                                                   .                                                                                                                                                                                                                       	    	      /                                                                                                                                                                                                           ,                                                                                                                                                                                                                             -                                                                                                                                                                                                                          .    	                                                                                                                                                                                                                         1                               	                                                                                                                                                                                     ,                                                                                                                                                                                                                             -                                                                                                                                 
                                                                                      -                                                                                                                                                                                                                 .                                                                                                                                                                                                                                ,                                                                                                                                                                                                                      /                                                                                                                                                                                                            /                  
                                                                                                                                                                                                      /                                                                                                                                                                                                                                       /                                                                                 
                                                                                                                                /                                                                                                                                                                                                                   .                                                                                                                                                                                                                  .                                                                                                                                                                                                                 -     	                        	                                                                                                                                                                                             -                                                                                                                                                                                                                    .                                                                                                                                                                                                                       /                                                                                                                                                                                                            0                                                                                                                                                          	                                                      0                                                                                                                                                                                                              
/                                                                                                                                                                                                   	             .                                                                                                                                                                                                                              /                                                                                                                                                                                                             .                                                                                                                                     	                                                        	                       
            1                                                                                                                                                                                                                       -                                                                                                                                                                                                                                .                                                                                    	                                                                                                                                     /                                	                                                                                                                                                                                    /                                                                                                                                                                                                                      0                                                                                                                                                                                                                    .                                                                                                                                                                                                                        ,                                                                                                                                                                                                                               .                                                                                                                                                                                                               
/                                                                                                                                                                                                                          .                                                                                                                                                                                                                 /                                                                                                                                                                                                                         
  /                                                                                                                                                                                                                          -                                                                                         	                                                                                                                                  .                                                                                                                                                                                                                       .                                                                                                                                                                                                                    
     	  1                
                                                                                                                                                                                                       .                                                                                                                                                                                                                 -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                         0                                                                                                                                                                                                                           -                                                                                                                                                                                                                    -                                                                                                                                                                                                                            -                                                                                                                                                                                                                                   0                          	                                                                                                                                                                                                .                                                                                                                                                                                                        	         -                                                                                                                                                                                                                   .                                                                                                                              	                                                                             	           .                                                                                                                                                                                                                      0                                                                                                                                                                                                                             .        
                                                                                                                                                                                                           ,                                                                                                                                                                                                         -    	                                                                                                                                                                                                                        0                                                                                                                                                                                                                    -                                                                                                                                                                                                                            0                                                                                                                                                                                                              .                                
                                                                                                                                                                                          .                                                                                                                                                                                                                        1                                                                                 	                                                                                                                               /                                 	                                                                                                                                                                                     -                                                                                                                                                                                                             0                                                                                                                                                                                                   2                                                                                                                                                                                                           1                                                                                                                                                                             	 	                                0                                                                                                                                                                                                                 .                                                                                                                                                                                                                           /                                                                                                                                                                                                        /                                                                                                                                                                                                                 .                	                                                                                                                                                                                                          -              	                                                                                                                                                                                                           
           0                                                                                                                                                                                                       
0                               
                                                                                                                                                                    	        - 	                                                                                                                                                                                                                        .                                                                                           	                                                                                                                              .                                                                                                                                  	                                                                                   .                            
                                                        
                                                                                                                  	              -                                                                                                                                                                                                                             0                                                                                                                                                                                                           
      .                                                                                                                                                                                                                        .                                                                                                                                                                                                                          	   -                	                                                                                                                                                                                                    -                                	 
                                                                                                                                                                              	              /      	                                                                                                                                                                                                                    .                                                                                                                                                                                                                            0                                                                                                                                                                                                               /                                                                                                                                                                                                                 ,                                                                                                                                                                                                                  	             -                                                                                                                                                                                                                         /                                                                                                                                                                                                                         /                                                                                  
                                                                                                                                    ,                                                                                                                                                                                                                        -                                                                                                                                                                                                          	            	        	0                                	                                                                                                                                                                                         .                                
                                                                                                                                                                               .       
                                                                                                                                                                                                                    .                                                                                                                                                                                                        
       .               
                                                                                                                                                                                                        .                                                                                                                                                                                                                     	          -                                                                                         	                                                                                                                               0                                                                                                                                                                                                           ,                	                                                                                                                                                                                                            -                                                                                                                                                                                                                    
   .              	                                                                                                                
                                                                                       3                                                                                                                                                                                                   
               -                            
                                                                                                                                                                                               /                                                                                                                                                                                                                       /                                                                                                                                                                                                              .                            	                                                                                                                                                                                       .                                                                                                                                                                                                                   /                                                                                                                                                                                                      .                                                                                                                                                                                     
                         2                                                                                                                                                                                                       /                                                                                                                                                                                                                   -                                                                                                                                                                                             	                                  /                                                                                                                                                                                                            	/                                                                                                                                                                                                         .                                                                                                                                                                                                                             /                                                                                                                                                                                                    	       
                    /                                                                                                                                                                                                          1                                                                                                                                                                                                               -    	   	                                                                                                                                                                                                                 /                                                                                                                                                                                                                 .                                                                                                                                                                                                                      -                                                                                    	                                                                                                                                  .   	                                                                                                                                                                                                                    .                                                                                                                                                                                     	                           	       /                                                                                                                                                                                                                  .                                                                                                                                                                                                                      	    .              
                                                                                                                                                                                                           ,                                                                                           
                                                                                                                                 ,      	   	                        
                                                                                                                                                                                              .                                                                                                                                                                                                                              .    
                                                                                                                                                                                                               .                                                                                                                                                                                                                       -                                                                                                                                                                                                            	             -                                                                                                                                                                                                                        /                                                                                                                                                                                                                 
           .                                                                                                                                                                                                                     -                                
                                                                                                                                                                                              -                                                                                                                                                                                                                          1                                                                                                                                                                                                                         -                                                                                             	                                                                                                                        /                                                                                                                                                                                                                       -                                                                                                                                                                                                       	           /                                                                                                                                                                                                                        -                                                                                                                                                                                                 
                      .                                                                                                                                                                                                                       /                                                                                                                                                                                                                    -                 
                                                                                                                                                                                                           .                                                                                                                                                                                                                      	    /                                                                                                                                                                                                               -                                                                                                                                                                                                           -                                                                                                                                                                                                                          -                                                                                             	                                                                                                                               	.                                                                                        	                                                                                                                              .                                  
 
                                                                                                                                                                                    .                                                                                                                                                                                                    	              /                                                                                                                                                                                                          1                                                                                                                                                                                                      0                                                                                                                                                                            	                                /                                                                                                                                                                                                          -                                                                                                                                                                                                                          	     .                                                                                                                                                                                                    .                                                                                                                                                                                                                    .                                                                                                                                                                                                                                0                                                                                                                                                                                                                   
      	     2                                                                                                                                                                                                       .                                                                                                                                                                                              	     	         -                	                                                                                                                                                                                                      1                                                                                                                                                                                                                         -                                                                                                                                       	                                                                                -                                                                                                                                                                                                                 -               	                                                                                                                                                                                                                    0                                                                                                                                                                                                                      ,                	                                                                                                                                                                                                               .                                                                                                                                                                                                                                .            	                                                                                                                                                                                                             ,                                                                                                                                                                                                               	              .                                                                                                                                                                                                                            -                                                                                                                                                                                                                   
         .                                                                                                                                                                                                    		               ,                                                                                                                                                                                                                     -                                                                                                                                                                                                                      0                                                                                                                                                                                                   	                
  .                                                                                                                                                                                                               	              0                                                                                                                                                                                                                          ,                                                                                                                                                                                                                            /                                                                                                                                                                                                                           	   /                                                                                                                                                                                                                           .                                                                                                                                                                                                                            -                                                                                                                                                                                                                          -                                                                                                                                                                                    	                   	       0                                                                                                                                                                                                              
/           	                                                                                                                                                                                                  	              
            /                                                                                                                                                                                                                   /                                                                                                                                                                                                                         	    /                                                                                                                                                                                                                    ,                                                                                      	                                                                                                                           "                 -  	                   	                                                                                                           	                                                                                          -                                                                                                                                                                                                                    -                              
                                                                                                                                                                                             3                                                                                                                                                                                                                 0                                                                                                                                                                                                                      .                                                                                    
                                                                                                                                      2                                                                                                                                                                                      
                            1                                                                                                                                                                                                .                                                                                                                                                                                                        -                                                                                                                                                                                                                       1                                                                                                                                                                                                     	           .                                                                                                                                                                                    	   	                           -   
                                                                                                                                                                                                                /                                                                                                                                                                                         
                                /                                                                                                                                                                                                                   /                                                                                                                                                                                                                                   /                                                                                                                                                                                                            -                                                                                                                                                                                        	            	            .                                                                                                                                                                                                                     -                                                                                                                                                                                                                      	      -                                                                                                                                                                                                                       /                                                                                       	                                                                                                                          -                                                                                                                                                                                                                               /                                                                                                                                                                                                                       -                                                                                                                                                                                                                      .                                                                                                                                                                                                                        .                                                                                                                                                                                                                           -                                                                                         	                                                                                                                                         .                                                                                                                                                                                                                  	                    /                                                                                                                                                                                                             -          	      	                                                                                                                                                                                                   	            -                                                                                                                                                                                                            ,                                                                                                                                                                                                                      -                                                                                                                                                                                                                       /                                                                                                                                                                                                                        
   .                                                                                                                                                                                                           .                                                                                                                                                                                                                               /                                                                                                                                                                                                               
 	    	.                                                                                                                                                                                                                            -                                                                                                                                                                                                                                 .                                                                                                                                                                                                                                .                                                                                                                                                                                                         	        0                                                                                                                                                                                                             /                                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                   /                                                                                                                                                                                                                              .                                                                                                                                                                                                                          ,                                                                                             	                                                                                                                                      -    
                                                                                                                                	                                                                                            -                                                                                                                                                                                                          ,                                 	                                                                                                                                                                                               /                                                                                                                                                                                                                .                                                                                                                                                                                                                            .        	                                                                            
                                                                                                                                       -                                                                                                                                                                                                                       0                                                                                                                                                                                                      0                                                                                                                                                                                                        ,             
                                                                                                               
                                                                                   .                                                                                                                                                                                                                     ,                                                                                                                                                                                                
                               ,                      
                                                                                                                                                                                           .                                                                                                                                                                               
                                 ,                                                                                                                                     
                                                                                            -                                                                                                                                                                                                                                   	      /                                                                                                                                                                                                       /                                                                                                                                                                                                                 -                                                                                                                                                                                                                   -                                                                                                                                                                                                                              .                                                                                                                                                                                                                           -                                                                                   
                                                                                                                                     ,   	   	                                                                                                                                                                                                                           0                                                                                                                                                                                                               /                                                                                                                                                                                                                           /                                                                                                                                                                                                                      
    .               
                                                                                                                        	                                                                                      ,                                                                                                                                                                                                              
	                -                                                                                                                                                                                                                                      .                                                                                                                                                                                                                              ,    	     
                                                                                                                                                                                                   	               -                                                                                                                                                                                                                 -           
     	                                                                                                                                                                                                      
             -                                                                                                                                                                                                               -                                                                                                                                                                                                                               1                                                                                                                                                                                                                 -    	                                                                                                                                                                                                                         .                                                                                                                                                                                                           	       
 /                                                                                                                                                                                                                      .                                    	                                                                                                                                                                                      .                                                                                    
                                                                                                                                    -                                                                                                                                                                                                                /                                                                                                                                                                                                               /           
          
                                                                                                                                                                                                  
                     0                                                                                   
                                                                                                                      1                                                                                                                                                                                                        
           
     -    
   	                                                                                                                                                                                                                 -                                                                                                                                                                                                                   #                /                                                                                                                                                                                                                           /                                                                                                                                                                                                                  ,    
                                                                                                                                                                                                                          0                                                                                        	                                                                                                                    1                                                                                                                                                                                                         0                                                                                                                                                                                                          .                                                                                                                                                                                                                 0                                                                                                                                                                                                    1                                                                                                                                                                                           	.                                                                                                                                                                                                              .                                                                                                                                                                                                                -                                                                                                                                                                                                                          3                                                                                                                                                                                                                  /                                                                                                                                                                                                                  -                                                                                                                                                                                                                       /          	                                                                                                                                                                                                   	                         0                                                                                                                                                                                                    	,                                                                                                                                                                                                                 	   -     	                                                                                                                                                                                                                -                                                                                                                                                                                                                              -                                                                                                                                                                                                                       -                                                                                                                                                                                                                       -                                                                                                                                                                                                                            ,                                                                                                                                                                                            	   	                            .                                                                                                                                                                                                                    -                                                                                                                                                                                                     
             ,                                                                                                                                                                                                                                    -                                                                                                                                                                                                                  
                ,                                                                                                                                                                                                                  	    ,                                                                                                                                                                                                                    	    	    /                                                                                                                                                                                                                          -                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                    -                                                                                                                                                                                                                              1                                                                                                                                                                                                                ,                                                                                                                                                                                                                                	     .                                                                                                                                                                                                                        .                                                                                                                                                                                                                         -                                                                                                                                                                                                                      -                                                                                                                                                                                                                         ,                      	                                                                                                                                                                                                        ,                                                                                                                                                                                                     	                            ,                     	                                                                                                                                                                                                             -                                                                                                                                                                                                                      -                                                                                                                                                                                                                                      -          	                                                                                                                                                                                                        ,                                                                                                                                                                                                                                 -                                                                                                                                                                                                                                    .                                                                                                                                                                                                                                 .                                                                                   	                                                                                                                           -                                  	                                                                                                                                                                                     ,                                                                                                	                                                                                                                                     	-                                                                                                                                                                                                                     
                 -                                                                                                                                                                                                                             ,                                  
                                                         
                                                                                                                                  -                                                                                                                                                                                                	                           -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                        -                                                                                                                                                                                                                         -                                                                                                                                                                                            
                            ,                                                                                                                                          
                                                                                       -                                                                                                                                                                                                                   ,                
                                                                                                                                                                                                               -                                                                                                                                                                                                                            .                                   
                                                                                                                                                                                	            -                                                                                                                                                                                                      	                  -                                                                                                                                                                                                               	           -                        	                                                                                                                                                                                                             ,     	                                                                                                                         	                                                                                             ,          
                          
                                                      	                                                                                                                                       ,                                                                                                                                                                                                                             -                                                                                                                                                                                                                                  -                                   	                                                                                                                                                                                                 ,                                                                                                                                                                                                                                 .                              	                                                                                                                                                                                                 -                                                                                                                                                                                                                    .                                                                                                                                                                                                                                -                	       	                                                                                                                                                                                                      .          
                                                                                                                                                                                               	              -                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                                  ,          !                                                                                                                                                                                                                             .                                                                                                                                                                                                                    ,                                                                                                                                                                                                    
                 	                  ,                                                                                                                                 	                                                                                               ,                                                                                                                                                                                                                          .                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                       -                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                          -                  

                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                            -     
                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                  	  .                  !                                                                                                                                                                                                                   .                                                                                                                                                                                                                                     ,                        	                                                                                                                                                                                                     ,                                                                                                                                                                                                        	   	 
                              .                                                                                                                                                                                                                        ,                                                                                                   		                                                                                                                                  
    ,                                    
                                                                                                                                                                                ,                                                                                                                                                                                                                                        -          	                                                                                                                                                                                                                              ,                                                                                                                                                                                                             
                                    ,                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                                   ,                                                                                                                                       	                                                                                                  ,                                                                                                                                                                                                                                               -                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                              	         .                                                                                                                                                                                                                      -                                                                                                                                                                                                                             ,           !                                                                                                                                                                                                                             ,                                                                                                                                                                                                                          $          -                
                                                                                                                                                                                                                 ,                                                                                                                                                                                                                            -                                                                                                                                                                                                                        -                                                                                                                                                                                                                                          -                                                                                                                                                                                                                                      -                                                                                                                                                                                                                                	     -                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                    -              
                                                                                                                                                                                                           ,                             	                                                                                                                                                                                           /                                                                                                                                                                                                                               ,                  	                                                                                                                                                                                                                   -               
                                                                                                                                                                                                          -                                  	                                                                                                                                                                                    ,                                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                .                                                                                                                                                                                                                     	      ,                                                                                                                                                                                                                               ,                                                                                                                                                                                                                     	      -                                                                                                                                                                                                                      
0                                                                                                                                                                                                                     -                                                                                                                                                                                                                                  ,               	       
                                                                                                                                                                                                             .                                                                                                                                                                                                	                          ,             

                                                                                                                      	                                                                                                ,                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                               -                                                                                                                                                                                                                             -                                                                                                                                                                                                                      -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                   -                                                                                                                                                                                                                           	        /                                                                                                                                                                                                                     ,                                                                                               	                                                                                                                               
-                                                                                                                                                                                                                                 .                                                                                                                                                                                                                              	-                                                                                                                                                                                                                                  -                                                                                                                                                                                                                     -                                                                                                                                                                                                                                     
.                                                                                                                                                                                                                           -                                                                                                                                     	                                                                                           ,                                                                                                                                                                                                                         	              -                  	                    
                                                                                                                                                                                              ,                                                                                                                                                                                                                                    -                  	                                                                                                                                                                                                     -                                                                                                                                                                                                                                        ,                  	                                                                                                                                                                                                             .                                                                                                                                                                                                                       .                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                      -                                                                                     
                                                                                                                                            ,                                                                                                                                                                                                                              	   	     ,                                                                                                                                                                                                                                    -                                                                                                                                                                                                                               ,                                     	                                                                                                                                                                                         /                                                                                                                                                                                                                             ,        	                                                                                                                      
                                                                                                    /                                                                                          	                                                                                                                            ,                                                                                                                                                                                                                              .         
          	                                                                                                                                                                                                             /                                                                                                                                                                                                                        ,                                                                                                                                      
                                                                            ,                                                                                                                                                                                                                             !         /                                                                                                                                                                                                                               0                                                                                                                                                                                                                        ,                                                                                                                                                                                                                              ,                                                                                                                                 	                                                                                   .                                                                                                                                                                                                                            ,                                                                                                                                                                                                                    /                                                                                                                                                                                        	                              -                                                                                                                                                                                                          -                                                                                                                                                                                                                	          -                                                                                                                                                                                                                                  -                                                                                                                                                                                                             
             -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                          ,                      	                                                                                                                                                                                                                ,                                                                                                                                                                                                                                ,       
                                                                                                                                                                                                                     .                                                                                                                                                                                                                             .                                                                                                                                                                                                                               -                                                                                                                                                                                                                  0                                                                                                                                                                                                                                     -                                                                                                                                                                                                              .                                                                                                                                                                                                                    -                                                                                                                                                                                                               
  
   ,                                                                                                                                                                                                       
                              	  	 1                                                                                                                                                                                                         	     .                                                                                                                                                                                                                          ,                                                                                                                                                                                                                       	                .                                                                                                                                                                                                  	                        
         ,                
                                                                                                                                                                                                	
            .                                                                                                                                                                                                                     ,                                                                                                                                                                                                                               -                                  
                                                                                                                                                                                          .           	                                                                                                                                                                                                                 -                                                                                                                                                                                                                              /                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                    -                                                                                                                                                                                                                               -        
     
                                                                                                                                                                                                                ,                                                                                                                                                                                                                                #       -                    
                                                                                                                                                                                                      ,                                       	                                                                                                                                                                                         .           	                                                                                                                    
                                                                                                 ,                                                                                              $                                                                                                                                    -                                                                                                                                                                                                           
    	          ,                 	                                                                                                                        
                                                                                          .                                                                                                                                                                                                          	             ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                                   !  	         -                      	              	                                                                                                                                                                                           -                                                                                                                                                                                                                            ,                                                                                                                                                                                                   	                 
                .                                                                                                                                                                                                                               ,                 	                                                                                                                                                                                                                  /                                	                                                                                                                                                                                      ,                                                                                                                                                                                                                                    -                                      G                                                                                                                                                                                                            ,                                       "                                                                                                                                                                                                    ,                                                                                                                                                                                                                                                  -                                                                                                                                                                                                               	           	    ,                                                                                                                                                                                                                       .                                                                                                                                                                                                                             .                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                    *            ,                )                                                                                                                                                                                                                           -                                                                                               	                                                                                                                                      -         
                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                          ,                                                                                             	                                                                                                                                            ,                                                                                            
                                                                                                                                  ,                                     $                                                                                                                                                                                                         -                                                                                                                                                                                                                            	        	  ,                                                                                                                                                                                                                                   	-                       
                                                                                                                   	                                                                                              ,                                                                                                                                    '                                                          
                                   -                                                                                                                                                                                                       
                                 -                         	                                                                                                                                                                                                                   -                                                                                                                                                                                                                                  .               
                                                                                                                                                                                                           -                                                                                                                                                                                                                                                  ,         	                                                                                                                                                                                                                               -                                                                                                                                                                                                                        !         -                                                                                                                                                                                                                                     ,                                                                                                 
                                                                                                                         
                ,                
                                                                                                                                                                                                              .                                                                                             	                                                                                                                                    ,                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                     -                                                                                                                                                                                                                              -                                                                                                                                                                                                              	           ,                                                                                                                                                                                                                                
,                                                                                                                                                                                                                       -                 	                                                                                                                                                                                                                         ,                	                                                                                                                                                                                                                 .                                                                                                                                                                                                                           -                                  	                                                                                                                                                                                       .                                                                                                                                                                                                                                     -                                                                                                                                                                                                                      .                                                                                                                                                                                                                     ,                                                                                                                                       	                                                                                           ,                                                                                                                                                                                                                                    .                                                                                                                                                                                                                          -                             
                                                                                                                                                                                      -                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                       
                            -                                                                                                                                                                                                  	                                   ,                                                                                                                                                                                                                                  !              -                !                                                                                                                                                                                                                           -                                                                                                                                                                                                                          
    ,                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                	     	     	 
  -                              	                                                                                                                                                                                                           -                                                                                            
                                                                                                                               ,                           	                                                                                                                                                                                            -                                                                                                                                                                                                                         	          	 
,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                              ,                                    	                                                                                                                                                                                      -                                                                                                                                                                                                                         
-                                                                                                                                                                                                                                    ,                                                                                                                                             #                                                                                                    -                                    
                                                                                                                                                        
                                      ,                                                                                                                                                                                                                                          .                	                                                                                                                                                                                                                      -                                                                                                                                                                                                                      
   -             	                                                                                                                                                                                                             ,                                                                                                                                                                                                                        	                        -         !                          
                                                                                                                                                                                              -                                                                                                                                                                                                                      -         	                                                                                                                                                                                                                     ,                                                                                               
                                                                                                                                     .         !       
       	                                                                                                                                                                                                                      .                                                                                                                                                                                                                                   ,                                   
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                   ,           
             
              
                                                                                                                                                                                           .                                                                                                                                                                                                                         -                                                                                                                                                                                                                      .                                                                                                                                                                                                                        
     	     ,                                                                                                                                                                                                                                   .                                                                                                                                                                                                                             ,                                                                                                                                                                                                                         .                                                                                                                                                                                                                                           -                                                                                                                                                                                                                                 /                                                                                                                                                                                                                              ,                                                                                                                                                                                                                               ,        	                                                                                                                                                                                                                  -                                                                                                                                                                                                                          .                                                                                                                                                                                                                     /                                                                                                                                                                                     
                      	         /                                                                                                                                                                                                                              .                                                                                                                                                                                                                        	     -             	    
     
                                                                                                                                                                                                               -                                                                                                                                                                                                                           	
              ,                   	                                                                                                                                                                                                                                 0                                                                                                                                                                                                                            .                                                                                                                                                                                                                               ,                                                                                                                                                                                                                   &              ,                                	                                                                                                                                                                                               -                                                                                                                                                                                                                          	       -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                        -                                                                                                    	                                                                                                                                      ,                                     
                                                                                                                                                                                            -                                                                                                                                                                                                                                         ,                                                                                                                                                                                                   
                      	       -                                                                                                                                                                                                                                   	     ,                       
                                                                                                                                                                         
                                    -                                                                                                                                                                                                                                 -                                                                                                                                                                                                   	                                    ,                 
                                                                                                                                                                                                                 ,                                                                                                                                                                                                                         -              	                                                                                                                                                                                                       ,                                                                                                                                                                                                                              ,                         	                                                                                                                                                                                                                       ,                                                                                                                                                                                                                   #      
          ,                                                                                                                                                                                                                                	     -                                                                                            
                                                                                                                                  -                                                                                                                               
                                                                                            -                                                                                          
                                                                                                                        
        	         /                                                                                                                                                                                                                                 0                                                                                                                                                                                                                         -                                                                                                                                                                                                           .               
                                                                                                                                                                                                        .                                                                                                                                                                                                                 -                              	                                                                                                                                                                         -         	                                                                                                                                                                                                         /                                                                                                                                                                                                                     	     	   /                                                                                                                                                                                              
            .                                                                                                                                                                                                                  0                                                                                                                                                                                                                     -           
                                                                                                                                                                                                        
           .                                                                                                                                                                                                                    2                                                                                                                                                                                                     
           /                           
                                                                                                                                                                            -                                                                                                                                                                                                      
                      .     	                        
                                                                                                                                                                                          .                                                                                                                                                                                                                   	,                                                                                                                                                                                                                               0                                                                                                                                                                                                        0                                                                                                                                                                                                               -                                                                                                                                                                                                                             0                                                                                                                                                                                                                    .                                                                                                                                                                                                                    /      	                                                                                                                                                                                                                 /                                                                                                                                                                                                                  /                                                                                                                                                                                                              .                                                                                                                                                                                                                 -                                                                                                                                                                                                                       1                                                                                                                                                                                                                  1                                                                                                                                                                                                                      3                                                                               	                                                                                                                               1                                                                                                                                                                                                                          1                                                                                                                                                                                                             /                                                                                                                                                                                                       -                                                                                                                                                                                	                            2                                                                                                                                                                                                        -                                                                                                                                                                                                                2                                                                                                                                                                                                     /                                                                                                                                                                                                        0                                                                                                                                                                                                                     /                                                                                                                                                                                                                          /                                                                                         	                                                                                                                    	          /                                                                                                                                                                                                                 0     	                                                                                                                                                                                                                     1                                                                                                                              	                                                                                     -                                                                                                                                                                                                                        -                                                                                                                                                                                                                            .                                                                                                                                                                                                                        -                                                                                                                                                                                                                                  0                                                                                                                                                                                             /                                                                                                                                                                                                                            .                                                                                                                                                                                                                .                                                                                          	                                                                                                                            -                                                                                                                                                                                                                   .                                                                                                                                                                                                            	         0                                                                                                                                                                                                               /                                                                                                                               	                                                                                .                                                                                                                                                                                                                    .          
                                                                                                                                                                                              	       	             -                                                                                                                                                                                                                    0                                                                                                                                                                                                    -                                                                                                                                                                                                             .                                                                                                                                                                                                      	                       .       
                                                                                                                                                                                                          -                                                                                                                                                                                                                 
.                                                                                     	                                                                                                                                       0                                                                                                                                 	                                                  	                               /                                                                                                                                                                                                           .                   	                                                                                                                                                                                                      .                                                                                                                                                                                                              	1                                                                                                                                                                                                           -                                                                                                                                                                                                                       0                                                                                                                                                                                                                           /                                                                                                                             
	                                                                                  0                                                                                                                                                                                                                  .                  
                                                                                                                                                                                                       /                                                                                                                                                                                                              1                                                                                                                                                                                                               /                                                                                    	                                                                                                                                         1                                                                                                                                                                                                          0                                                                                                                                                                               
                          /                                                                                                                                                                                         
                      /                                                                                                                                                                                      	                               -                                                                                                                                                                                                      .                                                                                                                                                                                                               0                                                                                                                                                                                                    /                                                                                                                                                                                                     -                                                                                                                                                                                                                      -                                                                                                                                                                                                                     /                                                                                                                                                                                                               		       1                                                                                                                                                                                                                   .                                                                                                                                                                                                                               /                 	                                                                                                                                                                                                ,                                                                                                                                                                                                                    ,       
                                                                             
                                                                                                                        	                -                                                                                                                                                                                                                         .                                                                                                                                                                                                                         /                                                                                                                                                                                                     /                                                                                                                                                                                                                         .                                                                                                                                                                                                                       1                                                                                                                                                                                                                -            
                                                                                                                                                                                                          /                                                                                                                                                                                                                       0                                                                                                                                                                                                        -                                                                                                                                                                                         	                             -                                                                                                                                                                                                                      -                                                                                                                                                                                                                           /                                                                                                                                                                                                                     0                                                                                                                                                                                                            0                                                                                                                                                                                                             1                                                                                                                                                                                              	                              
   -                                 	                                                                                                                                                                                      -       	                                                                                                                                                                                                           ,                                                                                                                                                                                                                       -                                                                                                                                                                                                                  /            
                                                                                                                                                                                                      .           
                                                                                                                                                                                                                   .                                                                                                                                                                                                  .                                                                                                                                                                                                 
        -                                                                                                                                                                                                                  .                                                                                                                                                                                                                    .                                                                                                                              
                                                                             /                                                                                                                                                                                                             -    	  	                                                                                                                                                                                                               1                                                                                    	                                                                                                                             	/                                                                                                                                                                                                               .                                                                                                                                                                                                                    2                                                                                                                                                                                                                    0                                                                                                                                                                                                        .                                                                                                                                                                                                          -                                                                                                                                      
                                                                                           /                                                                                                                                                                                                                -                                                                                                                                                                                                                 0                                                                                                                                                                                                    /                                                                                                                                                                                                            /                                                                                                                                                                                                                    /                                                                                                                                                                                                     	       	             0                                                                                                                                                                                                          	        0                                                                                                                                                                                                       .            	                                                                                                                                                                                                                    1                                                                                                                                                                                                              .                                                                                                                                                                                                                  -                             
                                                                                                                                                                                             0                                                                                                                                                                                                                           /                                                                                                                                                                                                                    	      .            	                                                                                                                                                                                       ,                                                                                                                                                                                                             	                 .                                                                                                                                                                                                                     /                                                                                                                                                                                                                       -                                                                                                                                                                                                    	                  .                                                                                                                                                                                                             "               .                                                                                                                                                                                                         0                                                                                                                                                                                                                 .          
     
                                                                                                                                                                                                 
             /                                                                                                                                                                                                         	             
   0                                                                                                                                                                                                            0                                                                                                                                                                                                                  ,     	                                                                                                                                                                                                      ,                                                                                                                                                                                                                                 ,                                   
                                                                                                                                                                                       -                                                                                                                                                                                                       /                                                                                              	                                                                                                                               -                                                                                                                                                                                                                  /                                                                                  	                                                                                                                              1                	                                                                                                                                                                                             -                                                                                                                                                                                                         
             0                                                                                                                                                                                                            ,                                                                                                                                                                                                                /                     
                                                                                                                                                                                                        .                                                                                                                                                                                                                /                                                                                                                                                                                                          /  
                                                                                                                                                                                                                        -                                                                                                                                                                                                            	          0                                                                                                                                                                                                                           -                          
                                                       	                                                                                                                                          0                                                                                          	                                                                                                                     /                                                                                                                                                                                                         	/                                                                                                                                                                                                         -                                                                                                                             
                                                                                      0                                                                                                                                                                                                            0                                                                                                                                                                                                      	           0                                                                                                                                                                                                                /                                                                                                                                                                                                   	         ,                                                                                                                            
                                                                                           /                                                                                                                                                                                                                        1                                                                                                                                                                                                                   /                                                                                                                                                                                                   -                    
                                                                                                                                                                                                          0                                                                                        	                                                                                                                       .                                                                                                                                  
                                                                               .                                                                                   	                                                                                                                        
                0                                                                                                                                                                                                           .                                                                                                                                                                                                                             -                                                                                                                                                                           	                               -                 	                                                                                                                                                                                                        -            
                                                                                                                     	                                                                                               .                         	                                                   
                                                                                                                              /                                                                                                                                                                                                                 .                                                                                                                                                                                                      	          
           -                                                                                                                                                                                                                       2                                                                                                                                                                                                   -                                                                                                                                                                                                                  .                                                                                                                                                                                                 	                    /                                                                                                                                                                                                                    .                                                                                                                                                                                                                     0                                                                                                                                                                                                                 /                                                                                                                                                                                                                           .                                                                                                                                                                                                                                  /                                                                                                                                                                                                                      /                                                                                                                                                                                                                   -                                                                                                                                                                                                       	      .                   	         	                                                                                                                                                                                             /                                                                                                                                                                                                                                       .                                                                                      	                                                                                                                                   0                                                                                                                                                                                                                 /   	                 	                                                                                                                                                                                                        -                                                                                                                                                                                                       	              -                    	                                                                                                                                                                                                     /                                                                                                                                                                                                            
            .   
                                       	                                                                                                                                                                             /                                                                                                                                                                                                                          2                                                                                                                                                                                                             /                                                                                   	                                                                                                                           .                                                                                                                                                                                                                     /                                                                                                                                                                                                             1                                                                                                                                                                                                     
-                                                                                                                                                                                                              2                                                                                                                                                                                                               -                                                                                                                                                                                        	                                /                                                                                                                                                                                                  	/                                                                                                                                                                                                               .                                                                                                                                                                                                                                   /                                                                                                                                                                                                           
               .                                                                                                                                                                                                         .                                                                                                                                                                                                          0                                                                                                                                                                                                                     /                                                                                                                                                                                                                          /                                                                                                                                                                                                                    -                                                                                                                                                                                                                            .                                                                                                                                                                                                         /                                                                                                                                                                                                   $                               0                                                                                                                                                                                                         -                                                                                                                                                                                                                            -                                                                                                                                         !                                                                                               0                                                                                                                                                                                                                        .           	                                                                                                                                                                                                              -                                                                                                                                                                                                                    .                                                                                                                                                                                                                         3                                                                                                                                                                                                    .        
                                                                                                                                                                                                                ,                                                                                                                                                                                                                       0                                                                                                                                                                                                                  .                                                                                                                                                                                                                     .                                                                                                                                                                                                            .                                                                                                                                                                                                                     .      
                                                                                                                                                                                                                                .                                                                                                                                                                                                            ,                                                                                        
                                                                                                                                        -         
                                                                                                                     	                                                                                       .                            	                                                                                                                                                                                                    1                                                                                                                                                                                                                                          0                                                                                                                                                                                                                         -                                                                                                                                                                                                            .   
              	                                                                                                                                                                                                       /                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                            .     
       	                  	                                                                                                                                                                                                  .                                                                                 	                                                                                                                         2                                                                                                                                                                                                                0                                                                                     
                                    	                                                                                   0                                                                                                                                                                                                                          .                                                                                                                                                                                                          /                                                                                                                                                                                                   
-                                                                                                                                                                                                               .                                                                                                                                                                                                       	             0                                                                                                                                                                                                                          /          	                                                                                                                                                                                              ,                                                                                                                                                                                                                       ,  	                                                                                                                                                                                                                                    /                                                                                                                                                                                                 
                      1                                                                                                                                                                                                     /                                                                                                                                                                                                                    .                                                                                                                                                                                                                           -                                                                                                                                                                                                                        -                                                                                                                                                                                                           	-                                                                                                                                                                                                                             0                                                                                                                                                                                                              /                                                                                                                                                                                                                                 ,                                                                                                                                                                                                       .                                                                                                                                                                                                 	                        -                                                                                                                                             )                                                                                    .                               
                                                                                                                                                                                    /      
                                                                                                                                                                                                      
                  0                                                                                                                                                                                                       
                        0                                                                                                                                                                                                                  -                                                                                                                                                                                                                  /                                                                                                                                                                                                                     /                                                                                                                                                                                                    
                    
       /                                                                                                                                                                                                           	        .                                                                                           	                                                                                                                         0        
                                                                                                                                                                                                    
,                                                                                                                                                                                                    	                       /                          "                                                                                                                                                                                                    ,                                      A                                                                                                                                                                                                     /        
                          
                                                                                                                                                                                             .                               
                                                                                                                                                     	                                 -                                                                                                                                                                                                                      ,             	                                                                                                                                                                                                          /                                                                                                                                                                                                    /                                                                                                                                                                                                               .                   	                                                                                                                                                                                       	             -                                                                                                                                                                                                                  $               ,                                                                                                                                   	                                                                                            .                                                                                                                                                                                                                        /                    
                                                                                                                                                                                                    .                                                                                                                                                                                                                 -                                                                                                                                                                                                                      /                                                                                                                                                                                                                     4                                                                                            	                                                                                                                     0                                                                                                                                                                                                         	/                                                                                                                                                                                                         	0                                                                                                                                                                                                                 	.                                                                                                                                                                                                                    .                                                                                                                                                                                           	                                  .                                                                                                                                                                                                          
/                                                                                                                                                                                                                    /                
                                                                                                           	                                                                                      .                                                                                                                                                                                                                                       2                                                                                                                                                                                                           .                                                                                                                                                                                                                   /     	     
                                                                                                                                                                                                               ,                                                                                                                                                                                                                       
        .                                                                                                                                                                                                                         -                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                   -                                                                                                                                                                                                $                               .              	                                                                                                                                                                                                  .                                                                                                                                                                                                                             ,                                                                                                                                     %                                                                                        /                                                                                                                                                                                                                .   
               	                                                                                                                                                                                                   .                                                                                                                                                                                                                                 /                                                                              	                                                                                                                         ,                                                                                                                                                                                      	                           -                                                                                                                                                                                                                 .                                                                                                                                                                                                                              /                                                                                                                                                                                                           /                                                                                                                                                                                                                       /        
                                                                                                                                                                                            -           
                                                                                                                                                                                               
       
                .                             #                                                                                                                                                                                   -                                      1                                                           
                                                                                                                                       -                                                                                                                                                                                                                    -                                                                                                                                                                                                                 .                                                                                                                                                                                                               .          
                                                                                                                                                                                                           -                                                                                                                                                                                                             .                                                                                                                                                                                                     
        ,                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                     /              	                                                                                                                                                                                                      .                                                                                                                                                                                                                 0    	                                                                                                                                                                                                                .                                                                                                                                                                                                                         -                                                                                             
                                                                                                                                0                                                                                                                                                                                                                        .                                                       	                                                                                                                                    
                          -                                                                                                                                                                                                      .                                                                                                                                                                                                                .                                                                                                                         
                                                                                           .                                                                                                                                                                                                                           -                                                                                                                                                                                                                           1                                                                                                                                                                                                     .                                                                                                                                 
                                                                                  -                                                                                                                                                                                                                 /          
                                                                                                                                                                                                                     /                                                                                                                                                                                                
-                                                                                                                                                                                                                -                                                                                                                                                                                                                          -                                                                                                                                                                                                                         -                                                                                                                                 	                                                                                      .                                                                                                                                                                                                                             -     
         
                  	                                                                                                                                                                                    -                                                                                                                                                                                                                          	          ,                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                      (         -                                                                                                                                                                                                                       /                                                                                                                                                                                                                    .    	    	          
                                                                                                                                                                                                               -                                                                                                                                                                                                                             
       0                   	                                                                                                                                                                                                          .                                                                                                                                                                                                      .                                                                                                                                                                                                                           -                                                                                                                                                                                                                                     2    	              
                                                                                                                                                                                     	          .                                                                                     	                                                                                                                        .                                                                                                                                                                                                                /                                                                                                                                                                                                                 '           /  	                                                                                                                                                                                                             -                                                                                                                                                                                                       	       /                                                                                                                                                                                                                    -                                                                                                                                
                                                     
                                 ,                                                                                                                                                                                                                .                                                                                                                                                                                                                                         -                                                                                                                                                                                                                          -                                                                                                                                                                                                          .          
                                                                                                                                                                                                             -                                                                                                                                                                                                                )                /                        	                                                                                                                                                                                      
                1                                                                                                                                                                                                             0                                                                                                                                                                                                                  ,                                                                                         	                                                                                                                             .                                 
                                                                                                                                                                                       -                                                                                                  	                                                                                                                               -                                                                                                                                                                                                                         /                                                                                                                                                                                                        .                                                                                                                                                                                  
                         /                                                                                                                                                                                                              1                                                                                                                                                                                                             -                                                                                                                                                                                                                               -                                                                                                                                                                               	                           3                                                                                                                                                                                           
                                 -                   	                                                                                                                                                                                                          /                                                                                                                                                                                                                                      -                                                                                                                                                                                                                      	         .                                                                                                                   
                                                                                        .       
                                                                                                                                                                                                       /                                                                                                                                                                                                               .                                                                                                                                                                                                                         ,                                 	                                                                                                                                                                                                   1       	                                                                                                                                                                                                        	-                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                   .                                                                                                                                                                                                                        #          /                                                                                                                                    '                                                                                         -                                                                                          
                                                                                                                               ,                                                                                                                                                                                                                    1                                                                                                                                                                                                                            /                                                                                                                                                                                                                    /                                                                                                                                                                                                                  .       
                                                                                                                                                                                               
              /                                                                                                                                                                                                      
               
  0                                                                                                                                                                                                               0                                                                                                                                                                                                                     .                                                                                                                                                                                                                  -                                                                                                                                                                                                                    -              1      
                                                                                                                                                                                                                 ,                                                                                                                                                                                  
                              	/                                                                                                                                                                                                                      .                                                                                                                                      	                                                                                       0                           	                                                                                                                                                                                       /                                                                                                                                                                                                                                 /                                                                                                                                                                                                                           0                                                                                                                                                                                                                .                                                                                                                                                                                                                  ,                                                                                                                                                                                                                 $               ,      
                                                                                     	                                                                                                                  
                 /                                                                                                                                                                                                                 /                                                                                                                                                                                                                 1                                                                                                                                                                                                           
-                                                                                                                                                                                                                             .                                                                                                  
                                                                                                                                  /                                                                                       
                                                                                                                              /                                                                                                                                                                                                              
.                                                                                                                             
                                                                             0                                                                                                                                                                                                                   
0                                                                                                                                                                                                /                                                                                                                                                                                                                    %          -                                                                                                                                                                                                                .                                                                                                                                                                                                                    ,   
                                                                                                                                                                                                                             .                                                                                                                                                                                                           	                        /                                                                                                                                                                                                             
                
   .                                                                                                                                                                                                                 /               	                                                                                                                                                                                               /                  	                                                                                                                                                                                                  -                                                                                                                                                                                                      
          -        
                          
                                                                                                                                                                                                /                 	                                                                                                                                                                                                       .                                                                                                                                                                                                                         
           -    	          		                                                                                                                                                                                                                  ,                                                                                                                                                                                                          
                            .                
                                                                                                                                                                                                              /                                                                               	                                                                                                                                  .                   	                                                                                                                                                                                                               -                                                                                                                                                                                                                                     /               
                                                                                                                                                                                                       -                                                                                                                                                                                                      -        	                                                                                                                                                                                                  	                -                                                                                                                                                                                                              
                 1     	                                                                                                                                                                                                                1                                                                                                                                                                                                                   /    	                                                                                                                                                                                                                  ,                                                                                                                                                                                                         !               /    
                                                                                                                                                                                                         .                                                                                                                                                                                 	                        .                                                                                                                                                                                                       -                  	                                                                                                                	                                                                                           ,                                                                                                                                                                                                                                /             	                                                                                                                                                                                                  	                       .                                                                                                                                                                                                                           
  -                                                                                                                                                                                                            -                                                                                                                                                                                                                        -                                                                                                                                                                                                               &             .                                                                                                                                                                                                                        0                           
                                                   	                                                                                                                                   /                                                                                                                                                                                                                  .                                                                                      
                                                                                                                             0                                   	                                                                                                                                                                                         -                                                                                                                                                                                                                                  /                                                                                                                                                                                      	                                      2                                                                                                                                                                                                        
/                                                                                                                                                                                                                -                                                                                                                                                                                                                .                                                                                                                                                                                                           -          	                                                                                                                                                                                                                      .                                                                                                                                                                                                              2                                                                                                                                                                                   	                             ,                                                                                                                                                                                                                            .                                                                                                                                                                                                        	                     0                                                                                                                                                                                                                       /       	                                                                                                                                                                                                  .                                                                                                                                                                                                              0                                                                                                                                                                                                              -                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                   .            
                                                                                                                                                                                                             -                                                                                                                                                                                           "                                  1                                                                                                                                                                                                                        ,                                                                                                                                  
                                                                                    -                                                                                                                                        '                                                        
                              .                                                                                                                                                                                                                     /                                                                                                                                                                                                         	             -                                                                                                                                                                                                                         
   ,                                                                                                                                                                                                               0                                                                                                                         
                                                                                 -                                                                                                                                                                                                                         	     /                                                                                                                                                                                                            	                 0                                                                                                                                                                                                                               -                                                                                               
                                                                                                                                /                                                                                                                                                                                                             /                                                                                                                                                                                                                      ,                                                                                                                                                                                                                           /                                                                                                                                                                                                                         ,                                                                                                                                                                                                                      -                                                                                                                                                                                                                  .                                                                                                                                                                                                                     -                                                                                                                                                                                                                                 .                                                                                                                                                                                                             /                                                                                                                                                                                                          .                                                                                                                                                                                                               ,        	                                                                                  
                                                                                                                            !                  .               	                                                                                                                                                                                                       0                                  	                                                                                                                                                                            -                                                                                                                                                                                                         .                                                                                    	                                                                                                                       
-                                                                                                                                                                                                                          .                                                                                                                                                                                                                     0                                                                                                                                                                                     
                               /                                                                                                                                                                                                                 /                                                                                                                                                                                                               .                                                                                                                          	                                                                                          3                                                                                                                                                                                                        ,                                                                                                                                                                                                                           .     	                                                                                                                                                                                                    1                                                                                                                                                                                   	                              -             	                                                                                                             
                                                                                      .                                                                                                                                                                                                               	                           /                                                                                                                                                                                                                 /                                                                                                                                                                                                      /                                                                                                                                                                                                         /                                                                                                                                                                                                                                -                                                                                                                                                                                                              /                                                                                                                                                                                                                   .                                                                                                                                                                                                                  -                                                                                               	                                                                                                                                	     ,                              
                                                                                                                                                                                            -                                                                                                                                                                                                              
           -                                                                                                                                                                                                                                 ,        
                                                                                                                                                                                                               
    -             	                                                                                                                     
                                                                                          -                                                                                                                                                                                                                                .                                                                                                                                                                                                                       -                                                                                                                                                                                                                           	   -          
                                                                                                                                                                                                                        ,         
                                                                                                                                                                                                                  .                                                                                                                                                                                                                     ,                                                                                                                                           	                                                                                       -        	  	                       
                                                                                                                                                                                              ,                                                                                                                                                                                                                   
    /                                                                                                                                                                                                                      -                                                                                                                                                                                                                                -                 
                                                                                                                                                                                                        -         	                                                                                                                                                                                                                      .                                                                                                                                                                                                                     ,                    
                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                       /                   
                                                                                                                                                                                                                  .                                                                                                                                                                                                              	               ,                                                                                                                                                                                                                                    -       	                                                                                                                                                                                                                                 /                                                                                                                                                                                                                               /                                                                                                                                                                                                                       -                   	                                                                                                                                                                                                               ,                                                                                                                                                                                                                             ,                                      -                                                                                                                                                                                           -                                                                                       
                                                                                                                                  ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                          	                       	    
    -                                                                                                                                                                                                 
                                 /                                                                                                                                                                                                                       ,                     /                                                                                                                                                                                                                           .          #           
                                                                                                                                                                                                                  .                                                                                                 
                                                                                                                        
            .                                                                                                                                                                                                                           
            -                                                                                                                                         	                                                                                                   ,                	                                                                                                                                                                                                  
                    ,            	                                                                                                                                                                                                                      ,                                                                                                                                                                                                                  #                ,                                                                                                                                      $	                                                                                            ,                                                                                                                                          8                                                                                               ,                                                                                                                                                                                                                           ,                                                                                                                                                                                                                 	                ,                                                                                                                                                                                                                          ,           ,               
                     	                                                                                                                                                                                        ,                                                                                                                                                                                                                               	   -                              	                                                                                                                                                                                                   -                                                                                                                                                                                                                            
      -              (                                                                                                                                                                                                                     ,                                                                                                                                                                                                                      (         .                 	                                                                                                                                                                                               -                                                                                                                                                                                                                         	                       ,                                                                                                                                                                                                                                       .                        	                                                                                                                                                                                                                     .                                                                                                                                                                                                                        -                                                                                                                                                                                                                                  -                                                                                      	                                                                                                                                      ,                   
                                                                                                                                                                                                             ,                               	                                                                                                                                                                                                 -                                                                                                                                                                                                                                    .                                                                                                                                                                                                                            ,                                 !                                                                                                                                                                                               .                                                                                                                                                                                                                 	     ,                                                                                                                                                                                                                               -          ,                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                       -     	                                                                                                                                                                                                                        	          ,                                                                                                  
                                                                                                                   	       '       	              ,                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                           
           -           
                                                                                
                                                                                                                                         ,                                                                                                      	                                                                                                                                             ,                                                                                                                                                                                                                                         	  ,                                  +                                                                                                                                                                                                             ,                                     -                                                                                                                                                                                                        ,                                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                              -                                                                                                                                           1                                                                                                   ,                     	                                                                                                                                                                                                                        ,                                                                                                                                                                                                  
                            '            ,                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                          
                   
     .                                                                                                                                                                                                                          -                                                                                                	                                                                                                                             %                    ,                %                                                                                                                         	                                                                                                   ,                                                                                                                                                                                                                                 	   	  	   .                    
                                                                                                                                                                                                          ,                                                                                                                                                                                                                                              2,                                                                                                                                                                                                                                              /                                                                                                 !                                                                                                                                      	.                                                                                                                                                                                                                            .        
                      
                                                                                                                                                                                      -                                   	                                                                                                                                                                                           -            
                                                                                                                                                                                                                 )          ,                
                                                                                                                                                                                                                   ,                                                                                                                                                                                                                       
              -            0                                                                                                                                                                                                                           -                                                                                                                                                                                                                                         -        	                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                    .       *                                                                                                                                                                                                                                    -                                                                                                                                                                                                                                    -                                                                                                                                                                                                                                         /                                                                                                                                                                                              	                      
   	      ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                               $            ,             	                                                                                                                                                                                                                ,                                     -                                                                                                                                                                                                   ,                                         -                                                                                                                                                                                                      -                               
                                                                                                                                                                                       ,                                                                                                                                                                                                                                ,                                                                                                                                                                                                          	                             	   /                                                                                                                                                                                                                          .                                                                                                                                                                                                                     
       .                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                  #                 -      
                                                                                                                                                                                                                   ,                                                                                                                                                                                                           
                                  /                                                                                                                                                                                                                          ,                                                                                                       
                                                                                                                            ,            
    ,                                                                                                     '                                                                                                                                           .                                                                                                                                                                                                                       - 
                                                                                                                                                                       
                                                    ,                                                                                                                                                                                                                 	                                ,                                                                                                                                                                                                              	                                      -                                                                                                                                                                                                                                .                                                                                                                                      	                                                                                         ,                                                                                                                                                                                                                                       	     ,                                                                                                                                                                                                                                ,                                           
                                                                                                                                                                                      
          -             
                                                                                                                                                                                                    -                                                                                                                                                                                                                       +                 /                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                          .                       
                                                                                                                                                                                             	         ,                                                                                                                                             -                                                                                           .                                                                                                                                                                                                                              /                                                                                                                                                                                                               .                                                                                                                                                                                                                      -                                                                                                                                                                                                                      -                                                                                                                                                                                                                          .                                     
                                                        
                                                                                                                                      .                                                                                                                                  	                                                                                     	,                                                                                                    	                                                                                                                          

             ,              	                                                                                                                                                                                                                -                                                                                                                                                                                                                                         .                                                                                                                                                                                                                      ,                                       
                                                            #                                                                                                                                       ,          
                       
                                                                                                                                                                                              .       
                                                                                                                                                                                                                       /      	                                                                                                                                                                                                         ,                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                              .                                                                                                                                                                                       	                              ,                                                                                              	                                                                                                                                   	   ,                              	                                                                                                                                                                                                -                                                                                                                                                                                                                                           ,                '                                                                                                                                                                                                                 -                                                                                                                                                                                                  
                               
      -                                                                                                                                                                                                                                      -                                                                                                                                                                                                          
           ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                   4                    .            "                                                                                                                                                                                                              -                                                                                                                                                                                                                                   ,                                  	                                                                                                                                                                                        ,                                                                                                     !                                                                                                                            
                 ,                                                                                                                                                                                                                                              -                                    $                                                                                                                                                                                                 -                                8                                                                                                                                                                                                     -                                                                                                                                                                                                               	             ,                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                     -                	                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                    (           ,         +                                                                                                                                                                                                                            -                                                                                                                                                                                                     	                                  ,                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                    	     -                                                                                                                                                                                                                        	               ,                                                                                           	                                                                                                                                     ,                                   	                                                                                                                                                                                                  ,                                                                                                                                                                                                                                   -                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                    ,                                     .  
                                                                                                                                                                                                 ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                        	                                   ,                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                           .                      
                                                                                                                                                                                                        ,                                                                                                                                                                                                         	                                        ,                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                           	              ,         
                                                                                                                                                                                                          .                                                                                                 &                                     
                                                                            	                ,                                                                                                                                                                                                                                    .                                                                                                                                                                                                                                       .                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                 
-                                                                                                                                                                                                                    
,                                     ;                                                                                                                                                                                                      ,                                  /                                                                                                                                                                                                        -                                                                                                                                                                                                                                  ,                                    '                                                                                                                                                                                                               -            	                        !                                                                                                                                                                                           -                                                                                                                                                                                                                                -                                                                                                                                                                                                                
     
           ,                                                                                                                                                                                                                                      .                                                                                                                                                                                                                                 ,             	                                                                                                                                                                                                                         ,                                                                                                  
                                                                                                                                       ,                                                                                                 	                                                                                                                                                ,                                                                                                   	                                                                                                                                      -                                                                                       	                                                                                                                                     ,                                                                                                                                             	                                                                                          ,                                                                                                                                                  	                                                           4                                     ,                                                                                                                                                                                                       +                                     ,                                                                                                                                                 E
                                                                                                    ,                                                                                                                                                                                                      .                                    ,                                    	                                                                                                                                                                                                               -                                                                                                                                                                                                    	                                    ,               
                                                                                                                                                                                                           /                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                                  -                                                                                                                                                                                                                               -             $                                                                                                                                                                                                              /                                                                                                                                           	                                                                                    .                                                                                                                                                                                                                              ,                                 	   
                                                                                                                                                                                                         -                                                                                                                                                                                                                           -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                     -                                                                                                                                                                                                                                 ,                                                                                                                                     
                                                                                                   ,                                                                                              	                                                                                                                                           .                 	                                                                                                                                                                                                     !                 -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                    .                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                	               .                                                                                                                                                                                                                            ,                                                                                                                                                                                                                   !                    ,                                     	                                                                                                 +                                                                                                 -                                                                                                                                                                                                                    	         -        	                            	                                                                                                                                                                                         ,                                                                                                                                  
                                                       
                                      ,       	                                                                                                                                                                                                                                   ,                                        "                                                                                                                                                                                             	       ,                         
                                                                                                                                                                                                                   ,                               	                                                                                                                                                                                    	,                   !                                                                                                                                                                                                                   
.                                                                                                                                                                                         	                                      ,                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                       ,           
       "                                                                                                                                                                                                                      -           	                                                                                                                                                                                                          "                -                      
                                                                                                                                                                                                        ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                  -                                                                                                    %                                                                                                                                      ,                                     0                                                                                                                                                                                                         ,                
       	                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                           ,                                                                                                 
                                      
                                                                                                ,                                                                                                     
                                                                                                                                           ,               $                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                            ,                                                                                                                                                   	                                                                                                ,                	                                                                                                                                                                                                                           -                                                                                                                                                                                                                                ,            '                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                   $               ,                        	                                                                     	                                                                                                                                             ,                
                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                      -                                                                                                  	                                                                                                                                ,         	                                                                                                                                                                                                                                         .                                                                                                                                                                                                                        ,                                                                                                                                                                                                                       ,                                                                                                                                                                                                                               -                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                     -             &      
                                                                                                                                                                                                                     ,                  	                                                                                                                                                                                                     %                -                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                       -                                                                                            	                                                                                                                                         -                                                                                                                                                                                                                                             -                                                                                                                                                                                                                            .                    	                                                                                                                   
                                                                          	             ,                                                                                                                                   
                                                                                      ,                                                                                                                                          
                                                                                           .                                                                                                                                                                                                                          ,      
                                                                                                                                                                                                                             ,                       
                                                                                                                                                                                                      /                                                                                                                                                                                                                        .                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                       -                                                                                                                                                                                                                                 .                                                                                                                                                                                                                                     /                                                                                                                                                                                                                    
          ,                                                                                                                                                                                                                              	,                                                                                                                                                                                                                                       /                                                                                                                                                                                                                      .                                                                                                                                                                                                                      ,             
                                                                                                                                                                                                                          ,                                                                                                       
                                                                                                                                    	     ,                                                                                                                                                                                                                                        -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                                 -                                                                                                                                                                                                                               ,                                                                                         	                                                                                                                               ,                                                                                                                                                                                                                                     -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                     /         	                                                                                                                                                                                                                         ,                
                                                                                                                                                                                                                               ,                                                                                                                                                                                                             .                                                                                                                                                                                                                             -                                                                                                                                                                                                                             -                                                                                          
                                                                                                                                    ,                                                                                                                              
                                                                                                 .                                                                                                                                                                                                            	                .                              
                                                                                                
                                                                                            ,                                                                                                                                                                                                                                ,                                   #                                                                                                                                                                                           -                                                                                                                                                                                                                             -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                -                                                                                                                                 
                                                                                         .                                                                                                                                                                                                                            0                                                                                                                                                                                                           -                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                         0               	                                                                                                                                                                                                             -                                                                                                                                                                                                                      -                               	  	                                                                                                                                                                                         ,                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                 -         
                         
                                                                                                                                                                                    .                                                                                                                                                                                                                              -                	                                                                            
                                                                                                                                      -                                                                                    
                                                                                                                                          .                                                                                                                                                                                                                                    -                                       
                                                                                                                                                                                     ,                                                                                                                                                                                                                           	           ,                                                                                                                                                                                                                                    -                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                  (            -         "                                                                                                                                                                                                                  ,                                                                                                                                                                                                                  
              -                                                                                                                                                                                                                                          -                                                                                                                                                                                                                   .                                  "                                                                                                                                                                                                   ,                                                                                                                                                                                                                         	     ,                                                                                                                                                                                                       !                                -                                                                                                                                                                                                                      /                                                                                                                                        #                                                                                                  ,                                                                                                                                                                                                                            *        0         !                                                                                                                                                                                                                      -                                     	                                                                                                                                                                               
               -                 
                                                                                                                       
                                                                                             ,                                                                                                                                                                                                                                -                  	                                                                                                                        	                                                                                            ,                                                                                                                                                                                                                                                 /              
                                                                                                                                                                                                                   ,                 
                                                                                                                                                                                                                   .            
                                                                                                                                                                                                              ,                                                                                                                                                                                                   	                              ,       
   	                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                            -                                                                                                                                                                                                                           -                                                                                                                                	                                                                                                ,                                                                                                                                                                                                                                         -                                                                                                                                                                                                                   !                    ,                                                                                                                                                                                                                               .                                                                                                                                                                                                                               ,                                                                                                                                                                                                                         /                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                              .                    	                                                                                                                                                                                                          .                                                                                                                                                                                                             	                ,                                                                                                                                                                                               	                             -                   	                                                                                                                                                                                                        .                
                                                                                                                                                                                                            -                                                                                                                                                                                                                                  .            	                                                                                 	                                        	                                                                                                      -                                                                                                                                                                                                             ,                                                                                                                                                                                                                                  .                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                    .       	                                                                                                                                                                                                  
    -           	    
                                                                                                                                                                                       	             ,                                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                      -                                                                                                                                                                                                                             -            
                                                                                                                                                                                                                        ,                                                                                               	                                                                                                                                      -                                   
                                                           	                                                                                                                                          ,                                                                                                                                                                                                               	         -                                                                                                                                                                                                                   ,                                                                                                                                                                                   	                             ,                                                                                                                                                                                                                                    .                                	                                                                                                                                                                                  -                                                                                                                                                                                                                -                                                                                                                                                                                                                                      ,        	                                                                                                                          
                                                                                               -                                                                                                                                                                                                                                  -                    	                                                                                                                                                                                                      .                                                                                                                                                                                                                	               -          !                                                                                                                                                                                                                       .                                                                                                                                                                                                                       -                                                                                                                                                                                                                                      /                                                                                                                                                                                                        
                -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                        	            .             
                                                                                                                                                                                                             ,                                                                                                                                                                                                                                           ,           	                      !                                                                                                                                                                                                        ,                                                                                               	                                                                                                                                           -              !                                                                                                                                                                                                                       ,       
                                                                                       	                                                                                                                                     .                                                                                                                                                                                                                                     	       ,                                                                                                                                        	                                                                                        -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                          
           -                                                                                                                                                                                                                                   +             ,                                                                                                                                                                                                                                              /                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                 ,                                  
                                                                                                                                                                                            ,                                                                                                                                                                                               
                  	      .                                                                                                                                                                                                                                ,                                                                                                                                                                                                           
   $                              ,                                                                                                                                                                                                                                        ,                               	                                                                                                                                                                                          .                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                   1   	      -                                                                                                                                                                                                          
                                      -                                                                                                                                                                                                                        .            -                                                                                                                                                                                                                                  -                                                                                                    
                                                                                                                                                ,                 &                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                           
          ,                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                       	           ,                                                                                                  '                                                                                                                                                  ,                                        4                                                                                                                                                                                                  .                                 	                                                                                                                                                                                    ,                                                                                                                                                                                                                                                
  ,                                                                                                                                                                                                               9                                   -                                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                                    ,                                                                                                                                                                                                    	                                        ,                                                                                                                                                                                                      	               .                                                                                                                                                                                                                           ,                                                                                                                                                                                                                              	       7              ,             (                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                   -                                                                                                                                                                                                                                    -                                                                                                                                                                                                                       "             
      ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                 .                                                                                                                                                                                                                     	        ,                                                                                                                                                                                                                      ,                                                                                                                                                                                                             .                                                                                                                                                                                                                       	     .                                                                                                                                                                                                                     .                              
                                                                                                                                                                                    -                                                                                                                                                                                                                           /                                                                                                                                                                                                                                   /                                                                                                                                                                                                                     0                                                                                                                                                                                     	                            .                                                                                                                                                                                                                  
           0                                                                                                                                                                                                                                   .                                                                                                                                                                                                              ,                                                                                                                                                                                                                            .                                                                                                                                                                                                                .                                                                                                                                                                                                                                .                                                                                                                                                                                                                   0                                                                                                                                                                                                      
     -     	                                                                                                                                                                                                                 /                                                                                                                                                                                                                - 	                                                                                                                                                                                                                      -                                                                                                                                                                                                                                      /                                                                                                                                                                                                               	-                                                                                                                                                                                                          .   	                                                                                                                                                                                                                      -                                                                                                                                                                                                                        "           -              
                                                                                                                                                                                                                -                                                                                                                                                                                                                          0                                                                                                                                                                                                                     1                                                                                                                                                                                                     .                                                                                                                                                                                                                     1                                                                                                                                                                                                               /                                                                                                                                                                                                          /                                                                                                                                                                                                   
-                                                                                                                                                                                                      .                	                                                                                                                                                                                                      .                                                                                                                                                                                 
                              .                                                                                                                                                                                                                         ,      	                         	                                                                                                                                                                                                      /                                                                                                                                                                                       	                                 0                                                                                                                                                                                                                  0                                                                                                                                                                                                                                         .                                                                                                                                                                                                           	/                                                                                                                                                                                                             -                                                                                                                                                                                                                           /                                                                                        
                                                                                                                                /                                                                                                                                                                                                                     /                                                                                          
                                                                                                                              ,   
  
   
      
      
                                                                                                                                                                                                          /                                                                                                                                                                                                              
        /                               	                                                                                                                                                          
                        /                  	                                                                                                                                                                                           	            	     -                                                                                                                                                                                                                           .                                                                                       	                                                                                                                              .                                                                                                                                                                                                                     /                                                                                                                                                                                                              
                          /                                                                                                                                                                                                                     0                                                                                                                                                                                                                  0        
                                                                                                                                                                                                           /                                                                                                                                                                                                                          0                                                                                                                                                                                                                  -                                                                                           
                                                                                                         	             .         	                                                                                                                                                                                                      ,                                                                                                                                                                                                                               .                             
                                                                                                                                                                                    0                                                                                                                                                                                                                   .                                                                                                                                                                                                                         .                                                                                                                                                                                                                 -                                                                                                                                                                                                                              .                                                                                                                                                                                                                                    -                
                                                                                                                                                                                                         -                                                                                                                                                                                                          .                    	                                                                                                                                                                                         -                                                                                                                                                                                                                       "              ,              #                                                                                                                                                                                                                     .                                                                                           
                                                                                                                  !                ,                                                                                                                                                                                                                    0                                                                                                                                                                                                        -                                     	                                                                                                                                                                                                 0                                                                                     	                                     
                                                                                                0                                                                                                                                                                                                                      .                                                                                                                                                                                                      -                                                                                                                                                                                                             .                                                                                                                                                                                                                   /                                                                                                                                                                                                            .                                                                                                                                                                                                                              ,      	                          	                                                                                                                                                                                                     /                                                                                                                                                                                                                         -                                                                                                                                                                                                                     .                                                                                                                                                                                                                     	                  -                                                                                                                                                                                                                 .                                                                                                                                                                                                                    .                                   
                                                                                                                                                                                                  0                                                                                                                                                                                                                             -                                                                                                                                                                                                            -                                                                                                                                                                                                                       -  
                  
                                                                                                                                                                                                   /                                                                                                                                                                                                                        /                                                                                                                                                                                                        0                                                                                                                                                                                                                           	  /                                                                                                                                                                                                                      .                                                                                     	                                                                                                                               /   	          
     
                                                                                                                                                                                                /                                                                                                                                                                                                                                    -                                                                                                                                                                                                                        .                                                                                                                                                                                                           .                                                                                                                                                                                                                  /                                                                                                                                                                                                                         /                                                                                                                                                                                                         	    /                                                                                                                                                                                                                  /                                                                                                                                                                                                                     .                                                                                                                                                                                                      	                        .                                                                                                                                                                                                                   0                                                                                                                                                                                                            	     ,                                                                                                                                                                                                                           -                                                                                                                                                                                                            -                                                                                                                                                                                                                                          .                                                                                                                                                                                                                   "                .                                   	                                                                                                                                                                                          ,                                                                                                                                                                                                                 .                                                                                                                                                                                                                       .                                                                                                                                                                                                                        #            ,                                                                                                                                                                                                                             -                                                                                            	                                                                                                                               -                     	                                                                                                                                                                                                  .                                                                                    
                                                                                                                          /                                    	                                                                                                                                                                                                ,                                                                                        	                                                                                                                                  .                                                                                                                                                                                                                                     0                                                                                                                                                                                                1                                                                                                                                                                                 	                           /                                                                                                                                                                                                                -                                                                                                                                                                                                             .                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                 /                                                                                                                                                                                                                       -           
                                                                                                                                                                                                          -                                                                                                                                                                                                                                        ,       	                                                                                                                                                                                                    ,                                                                                                                                                                                                     	               -                                                                                                                                                                                                                                  /                      	                                                                                                                                                                                                         ,                                                                                                                                                                                                                   ,                                                                                                                                                                                                                  ,  
                                                                                                                                                                                                                        .                                                                                                                                                                                                	                           	         -               
                                                                                                                                                                                                                    /                                                                                                                                                                                                                       -                                                                                                                                                                                                                        ,                                  
                                                      	                                                                                                                                   -      	   
                                                                                                                                                                                                                     ,                                                                                                                                                                                                         	                     .                                                                                                                                                                                                                          ,                                                                                                                                                                                                                 /         
      
                                                                                                                                                                                                                 /                                                                                                                                                                                                      
                	1                                                                                                                                                                                                                /                                                                                                                                                                                                                 ,                                                                                                                                                                                                                          /                                                                                                                                                                                                                            /                                                                                                                                                                                                                           .                                                                                                                                                                                                              -                                                                                                                                                                                                                              .                                                                                                                                                                                  
                                    -                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                     .                                                                                                                                                                                                                   -                                                                                                                                                                                                                .                                                                                                                                                                                                                        .                  	                                                                                                                                                                                                                   .                	                                                                                                                                                                                                -                                                                                                                                                                                                             /                                                                                                                                                                                                                /                                                                                                                                                                                                                   	.                                                                                                                                                                                                                 .                                                                                          	                                                                                                                        -                                                                                                                                                                                             	                              /                                                                                                                                                                                	                           1                                                                                                                                                                                                          
.                                                                                                                                                                                                               .                                                                                                                                                                                                                  .          	           	                                                                                                                                                                                                                -                                                                                                                                                                                                               .                                                                                                                                                                                                                     -                                                                                                                                                                                                                          -         
                                                                                                                                                                                                                            0                                                                                                                                                                                                         .                                                                                                                                                                                                            ,                                  	                                                                                                                                                                                       /                                                                                                                                                                                                                 /                	                                                                                                                      
                                                                                     /                                                                                                                                                                                                                       .                  	                          	                                                                                                                                                                           	/                                                                                                                                                                                             	                                ,                     	                                                                                                                                                                                                       -                                                                                                                                                                                                                  	                  .                                                                                                                               		                                                                                        /                                                                                                                                                                                                                     ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                     	   -             	                                                                                                                                                                                                                   .                                                                                                                                                                                                           ,       
                                                                                                                                                                                                                       .                                                                                                                                                                                                       
        /          
                                                                                                                                                                                                     .                                                                                                                                                                                                                   -     	                                                                                                                                                                                                                         .                                                                                                                                                                                                           
      
        	/      	                                                                                                                                                                                                 
                   /                                                                                                                                                                                                                .   
                                                                                                                                                                                                                  -                                                                                                                                
                                                                                       ,           	                  	                                                                                                                                                                                      /                                                                                                                                                                                                                                     -                                                                                                                                                                                                                 
  /                                                                                                                                                                                                                     .                 	                                                                                                                                                                                                    /                     
                                                                                                                                                                                                             -                                                                                                                                                                                                                      /                                 	                                                      
                                                                                                                        -      
                                                                                                                                                                                                                  0                                                                                                                                                                                                                      .                                                                                                                                                                                                                        .                                                                                               
                                                                                                                             .                                                                                                                                                                                                                                0                                                                                                                                                                                                          1                                                                                                                                                                                                      0                                                                                                                                                                                               0                                                                                                                                                                                                                   .                                                                                                                                                                                                                             -                                                                                                                                                                                            	                        
      .                                                                                                                                                                                            	                      	         -                                                                                                                                                                                                                                 .                                                                                                                                                                                                                                     .        	                                                                                                                                                                                                            0                                                                                                                                                                                                             ,                                  
                                                                                                                                                                                      /                                                                                                                                                                                                              ,                                                                                                                                                                                                                            ,                                                                                                                                                                                                                          -                                                                                                                                                                                                                 -                                                                                                                                                                                            
                              
      ,              	                                                                                                                                                                                                       .                                                                                                                                                                                                                              /            
                                                                                                                  	                                                                                          ,                                                                                                                                                                                                                         .                          	                                                                                                                                                                                               -                                                                                                                                                                                                               	                  .                                                                                     
                                                                                                                    	                ,                                                                                                                                                                                                           -                                                                                                                                                                                                                  .                                                                                                                                                                                                                           -                                                                                                                                                                                                              /                                                                                                                                                                                                                          -              
                                                                                                                                                                                                           .                                                                                                                                                                                                                         1                                                                                                                                                                                                                           /                                                                                                                                                                                                                    ,                                                                                                                                                                                                                       -                                                                                                                                                                                                                            2                                                                                                                                                                                                               -              
                                                                                                                                                                                                                     -                                                                                                                                                                                                                           .                                                                                                                                                                                                                    -  	                                                                                                                                                                                                                  /                                                                                                                                                                                                                                    .                                                                                                                                                                                                            .                             	                                                                                                                                                                                       -                                                                                                                                                                                                                      3                                                                                                                                                                                                             .                         
                                                                                                                                                                                            -                                                                                                                                                                                                                              /                                                                                                                                                                                                                       /                                                                                                                                                                                                 	/                                                                                                                                                                                                            .                                                                                                                                                                                  
                            1                                                                                                                                                                                                                    .                                                                                                                                                                                                                          .    
      	                                                                                                                                                                                                           /                                                                                                                                                                                            !                        	          .          
                                                                                                              
                                                                                        -                                                                                                                                                                                                                       .                                                                                                                                                                                                                     1                                  	                                                                                                                                                                                    -    	                                                                                                                                                                                                                 1                                                                                                                                                                                                     	             	-               
                                                                                                                                                                                                             ,                                                                                                                                                                                                                         .                                                                                                                                                                                                                      ,                                                                                                                                                                                                  	  #                               -                                                                                                                                                                            	                                  ,                                                                                                                                                                                                                                          ,              	                                                                                                                      
                                                                                         -                                                                                                                                                                                                                                -                                                                                                                                                                                                                              .                                                                                                                                                                                                                   	 1            	                                                                                                                                                                                         	                .                                                                                                                                 	                                                                               /                                                                                                                                                                                                                               -                                                                                                                                                                                                                  
      /                                                                                                                                                                                                                   ,                                                                                  	                                                                                                                                          /                                                                                                                                                                                                                       -                                                                                                                                                                                                                                  !       -                                                                                                                                                                                                                      /                                                                                                                                                                                                               ,      	                                                                                	 	                                                                                                                                             -                                                                                                                                	                                                                                        -              	                 	                                                                                                                                                                                                 /                                                                                                                                                                                                                        
             1                                                                                                                                                                                                           0                                                                                                                                                                                                             .              
                                                                                                                                                                                                               /         
                                                                                                                                                                                                                 .                                                                                                                                                                                                                  1                                                                                                                                                                                               
            -                    	            	                                                                                                                                                                                         -                                                                                                                                                                                                                      	 /                                                                                                                                                                                                                  /                                    	                                                                                                                                                                               /                                                                                                                                                                                                                           0                                                                                                                                                                                                                 /                                                                                                                                                                             
                           -                                                                                                                                                                                      	                               	/                                                                                                                                                                                    	                          -                                                                                                                                                                                                                                  1                                                                                                                                                                                                            -                                                                                                                                                                                                                   0                                                                                                                                                                                                                        ,                                                                                                                                                                                                   	                         .                                                                                                                                                                                                    0                                                                                                                                                                                                            -                                                                                                                                                                                                                     /                                                                                                	                                                                                                                           -             

                                                                                                                                                                                                         .                                                                                                                                                                                                                     -                                                                                                                                                                                                                                     .                                                                                                                                                                                            	  &                                      /                                                                                                                                                                                                           .                                                                                                                                                                                                                    -                                                                                                                                                                                              	                          .                                                                                 
 
                                                                                                                                  0            	                                                                                                                                                                                                   1                                                                                                                                                                                                                            
      0                                                                                                                                                                                                                       .                                                                                                                                                                                                         -                                                                                                                                                                                                                       .            	                                                                                                                                                                                                                          0                                                                                                                                                                                                                   /                                                                                    
                                                                                                                               /                                                                                                                                                                                                             /                                                                                                                                                                                                                            /                                                                                                                                                                                                                 -                                                                                                                                                                                                              -                                                                                
                                                                                                                                       -                                                                                                                                                                                                                   -                   	                                                                                                                                                                                                         0                                                                                                                                                                                                                           -                                                                                                                                                                                                             /                                                                                                                                                                                                	         .              	                                                                                                                                                                                                        /                                                                                                                                                                                                                     
    .                                                                                                                                                                                                                   ,                                                                                                                                                                                                       .                                                                                                                                                                                                                        .                                                                                     	                                                                                                                  	              	2                                                                                                                                                                                                                
-                                                                                                                                                                                                                       0                                                                                                                                                                                                                     1                                                                                                                                                                                                       1                                                                                                                                                                                                                 /                                                                                                                                                                                                                    0                                                                                                                                                                                                                      ,                                                                                                                                                                                              	                               .                                                                                                                                                                                                         /                                                                                                                                                                                                      -                                                                                                                                                                                                                      .             
      	                                                                                                                                                                                                              2                                                                                                                                                                                                             /                                                                                                                                                                                                             /                   	                                                                                                                                                                                                    /                                                                                                                                                                                                         
           1               
                                                                                                                                                                                                   -                                                                                       
                                                                                                                                    ,                                                                                                                                                                                                                               -                                                                                                                                                                                                  "                          
       .                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                  -                                                                                       	                                                                                                                                 -                                                                                                                                                                                                                              /                                                                                                                                                                                               	                	 ,                 
                                                                                                                                                                                                       -                                                                                                                                                                                       	                               -                                                                                                                                                                                                                             /                                                                                                                                                                                                                        0                 
                                                                                                                                                                                                     -                                                                                      	                                                                                                                                  -                             	                                                                                                                                                                                      ,                                                                                                                                                                                                                                  .      
                        
                                                                                                                                                                                          /                                                                                                                                                                                                               -                          
  
                                                                                                                                                                                    ,                                                                                                                            	                                                                                      ,                          
                                                    	                                                                                                                                         /                	                                                                                                                                                                                                       
      .                                                                                                                                                                                                                    /                                                                                                                                                                                                              -   	                                                                                                                                                                                                                         /         
                                                                                                                                                                                                                 .                                                                                                                                                                                                                  .                                                                                                                                                                                                                    .                                                                                                                                                                                                                           /                                                                                                                                                                                                                   /                                                                                                                                                                                                                  2                                                                                     
                                                                                                                         /                                                                                                                                                                                                                     2                                                                                                                                                                                    	                       	0                                                                                                                                                                                                     .                                                                                                                                                                                   	                              0                                                                                                                                                                                                                  	-                                                                                                                                                                                                                              .                                                                                                                                                                                                  /                                                                                                                                                                                                              -                                                                                                                                                                                                             1                                                                                                                                                                                                               
              	    2                                                                                                                                                                                                                2                                                                                                                                                                                                                 .                                                                                                                                                                                                                          .                                                                                                                                                                                                         
              .              
                                                                                                                      	                                                                                    -                                                                                                                                                                                                                          -                                                                                                                                                                                                                               -                                                                                                                                                                                                                  -           	                                                                                                                                                                                               /                                                                                                                                                                                                                          .                                                                                                                              
                                                                                           /                                                                                                                                                                                                                                .       
                                                                                                                                                                                                                       /                                                                                                                                                                                                               -                                                                                                                                                                                                                              2                                                                                                                                                                                                           .                                                                                                                                                                                                                       
      
     2                                                                                                                                                                                                            .                                                                                                                                                                                                               	              
   /                                                                                                                                                                                                       	               -                                                                                                                                                                                                                       1                                                                                                                                                                                                             	0                             
                                                                                                                                                                                 	          -                                                                                                                                                                                                                         -                                                                                                                                                                                                                       .                                                                                                                                                                                                               /   
                                                                                                                                                                                                          .                	                                                                                                                                                                                                                             /                                                                                                                                                                                                               /                                                                                                                                                                                                                          -            
                                                                                                                                                                                                             -                                                                                                                                                                                                                                   -  	                                                                                                                                                                                                                    1                                                                                                                                                                                                                      -      
                                                                                                                                                                                                             5                                                                                                                                                                                                      1                                                                                                                                                                                                                2                                                                            	                                                                                                                                  0                                                                                                                                                                                                          	         2                                                                                                                                                                                                          	1                                                                                                                                                                                                      	-                                                                                                                                                                                                             0                                                                                                                                                                                                                 	/                                                                                                                                                                                                                               .         	                                                                                                                                                                                            -                                                                                                                                                                                                                  -                                                                                                                                                                                                                     .              
                                                                                                                                                                                                	              
             0                                                                                                                                                                                                         -         	                                                                                                                                                                                                         /                                
                                                                                                                                                                                       .                                                                                                                                                                                                                               -                                                                                                                                    		                                                                             0                                                                                                                                                                                                                
              0       	         	                                                                                                                                                                                                           .                                                                                                                                                                                                                          -                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                        .                                                                                                                                                                                                                      1                                                                                        
                                                                                                                        /                   	                                                                                                                                                                                                        .                                                                                                                                                                                                                             0                                                                                                                                                                                                                   .                                                                                                                                                                                                          
         .                                                                                                                                                                                                                          /                                                                                                                                                                                                                               .                  
                                                                                                                                                                                                 0                                                                                                                                                                                                         1                                                                                                                                                                                                                  .                                                                                                                                                                                                                                   .                            
                                                                                                                                                                                          0                                                                                                                                                                                                               .                                   	                                                                                                                                                                                        -           
                                                                                                                                                                                                       
           0                                                                                                                                                                                                                      /                                                                                                                                                                                                              
        .                                                                                                                                                                                                                   -             	                                                                                                                                                                                                 /                                                                                                                                                                                                                                 0                                                                                                                                                                                                         
            .                                                                                                                          	                                                                                        .                                                                             	                                                                                                                             .      
                                                                                                                                                                                                                           .                                                                                                                                                                                                                ,                                    
                                                                                                                                                                                            -                          
                                                                                                                                                                                            3                                                                                                                                                                                                                 .                                                                                                                                                                                    
                            0                                                                                                                                                                                                                              -                                                                                                                                                                                          	                                     .                                                                                                                                                                                                            .                                                                                                                                                                                                                /          
                                                                                                                                                                                                        0                                                                                                                           	                                                                                 /                                                                                                                                                                                                                         .                                                                                                                                                                                                                          	     .                                                                                                                                                                                                  
            /                                                                                                                                                                                                           -  
                                                                                                                                                                                                                      2                 
                                                                                                                                                                                                /                                                                                                                                                                                                                       ,      
                        	                                                         	                                                                                                                                              .                                                                                                                                                                                                                  .                                                                                                                                                                                                                                 .                
                                                                                                                  	                                                                                    /                                                                                                                                                                                                     	                 .                                                                                                                                                                                                                    /                                                                                         	                                                                                                                      .                    	                                                                                                                                                                                                          -                                                                                                                                                                                                                                    /                                                                                                                                                                                                          
       -                                                                                                                                                                                                                  -                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                     .          
                                                                                                                                                                                                             1                                                                                                                                                                                                          -                                                                                                                                                                                                                   .                                                                                                                                                                                                              	              .                                
                                                                                                                                                                                     /                                                                                                                                                                                                                -                                                                                          	
                                                                                                                                   -             
                                                                                                                                                                                                         /                                                                                                                                                                                                                            /                                                                                                                                                                                                                                      1                                                                                                                                                                                                                      0                                                                                                                    	                                                                                     .                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                   0                                                                                                                                                                                                    -                                                                                                                                                                                                             -   
                           	               	                                                                                                                                                                              /                                                                                       	                                                                                                                                  -                                                                                              	                                                                                                                                     .  
               	                                                                                                                                                                                                          /                                                                                                                                                                                                   .                                                                                                                                                                                                               	/                                                                                                                                                                                                                 -                                                                                                                                                                                                                              0                                                                                                                                                                                                         -                                                                                                                                                                                                       -                                                                                                                                                                                                       /                                                                                                                                                                                                            /                                                                                                                                                                                                                      /                                                                                                                                                                                                                              1                                                                                                                                                                                                                       /                                                                                                                                                                                                             -                                                                                                                                                                                                                       0                                                                                                                                                                                                                    -                                                                                                                                                                                                                         -                                                                                                                                                                                                                               0                                                                                                                                                                                                                          -                                                                                                                                                                                        
                                   0           		                                                                                                              
                                                                                      .                                                                                                                                                                                                                        	              -                                                                                                                               	                                                                                       2                                                                                       	                                                                                                                          ,          
     	       
                                                                                                                                                                                                               -                                                                                                                                                                                                            
/                                                                                                                                                                                                              .                                                                                                                           
                                                                              -                                                                                                                                                                                                                          .                                                                                                                                                                                                          .                                                                                                                                                                                                                          .                                                                                                                                                                                                                           -  	                      	                                                                                                                                                                                            /                                                                                                                                                                                                          	  /                                                                                                                                                                                                           	                  .                                                                                                                                                                                                                    -            	                                                                                                                                                                                                                              .                                                                                                                               	                                                                             
          /                                                                                                                                                                                                                     -                                                                                                                                                                                                     	               
     0                                                                                                                                                                                                           	.                                                                                                                                                                                                         ,              	                                                                                                                                                                                                                     /                                                                                                                                                                                                                         1                                                                                                                                                                                                            .                                                                                                                                                                                                 	              0                                                                                                                                                                                                                             .                                  
                                                                                                                                                                                         0                                 	                                                                                                                                                                                             ,            	                                                                        
                                                                                                                                               0                                                                                                                                                                                                             .                                                                                                                                      	                                                     
                        1                                                                                                                                                                                                                      ,                                                                                                                                                                                              
                                   4                                                                                                                                                                                                            -                                                                                                                                                                                                         /                              
                                                                                                                                                                                  .                                                                                                                            
                                                                                 .              
                                                                                                                    
                                                                                         -                                                                                                                                                                                                                         /                                                                                        
                                                                                                                            2                                                                                                                                                                                                              /                                                                                                                                                                                                                          0                                                                                                                                                                                                              ,                                                                                                                                       	                                                                    	          -                                                                                                                                                                                                                               .                                                                                                                              	                                                                                                 -                                                                                                                                                                                           ,                            	        ,                                                                                                                                                                                                                  -                                                                                                                                                                                                                     /             	                                                                                                                                                                                                                         -                                                                                                                                                                                                                             -                                                                                                                                                                                                                                    -                                                                                                                                                                                                                                /                                                                                                                                                                                                                     .                                                                                                                                                                                                   ,                                                                                                                                                                                                                   	         .                                                                                                                                                                                                                     	0         
                                                                                                                                                                                                             .                                                                                                                           	                                                                                        -                                                                                                                                                                                                                  /                                                                                                                                                                                                          0                                                                                                                                                                                                                     -                                                                                                                                                                                                             .                                                                                                                                                                                                                             .                                                                                                                                                                                                                ,                                                                                                                                                                                                                     /                    
                                                                                                                                                                                                          /                                                                                                                                                                                                                     0                                                                                                                                                                                                                0                                                                                                                                                                                                                        .                                                                                                                                                                                                                 -                       	                                                                                                         	                                                                                                .                                                                                          
                                                                                                                     "                 -                    	          
                                                                                                                                                                                                 -                                                                                                                                                                                                                              .                                                                                                                                                                                                                             -                                                                                                                                                                                                                          /                                                                                         	                                                                                                                              ,                                                                                                                                  
                                                                               /                                                                                                                                                                                                         .                                                                                                                                                                                    	                                    -                                                                                                                                                                                                              .                                                                                                                                                                                                                  -                                                                                                                                                                                                           	-                                                                                                                                                                                          
                            
  -                                                                                                                                                                                                                                        /                                                                                                                                                                                                                    
   3                                                                                                                                                                                                           /                                                                                                                                                                                                            .                                  	                                                                                                                                                                                      0                                                                                                                                                                                                                     -                                                                                                                                                                                                                           .                                                                                                                                                                                                                              /                                                                                                                                                                                                            .                                                                                                                                                                                             ,                                   ,             
                                                                                                                                                                                                           -                                                                                                                                                                                                                    	   
     	 -             (      	                                                                                                                      	                                                                                                     1                                                                                                                                                                                                                              -                                                                                                                                                                                                                               -                                                                                                                                                                                                                 	        	   1                                                                                                                                                                                                                  /                                                                                                                                                                                                            -                                                                                                                                                                                                                      .                                                                                                                                                                                                                  /                                                                                                                                                                                                               -                                                                                                                                                                                                             -                                                                                                                                                                                                                           /                                                                                                                                                                                                                /                                                                                                                                                                                                                             .                                                                                                                                                                                                                  1                                                                                                                                                                                                                       1                                                                                                                                                                                                                  /                                                                                                                                                                                                                    /                      
                                                                                                                                                                                                             ,                                                                                                                                                                                                              	               /                                                                                                                                                                                                                 -                    	                                                                                                                                                                                                        0                                                                                                                                                                                                
                	    -                                                                                                                                                                                                                         
.                                                                                                                                                                                                                       .       	                        	                                                                                                                                                                                           -                                                                                                                                                                                                                                 /                                                                                                                                                                                                                         -                                                                                                                                                                                                                    ,                                                                                                                                                                                                                     -                                                                                                                                     	                                                     	                          -                                                                                                                                                                                                           -                                                                                                                                                                                     	                                    /                                                                                                                                                                                                          /                                                                                                                                                                                                             	      
  0                                                                                                                                                                                                       
.                                                                                                                                                                                                               .                                                                                                                                                                                                                                   .                                                                                                                                                                                                                       .                                                                                                                                                                                                            /                                                                                                                                                                                                                      ,                                                                                                                                                                                                                             1                                                                                               	                                                                                                                     1                                                                                                                                     	                                                                              -                                                                                                                                                                                                                                   /                                                                                                                                                                                                        /                                                                                                                                                                                                                             -                                                                                                                                                                                                                  2                                                                                                                                                                                                            .       
           
                                                                                                                                                                                                     	             1                                                                                                                                                                                                                       - 	                                                                                                                                                                                                     
                /                                                                                                                                                                                                    	              4                	                                                                                                                                                                                                    	2                                                                                                                                                                                                      	-                                                                                                                                                                                                                           1                                                                                                                                                                                                  
          	0    
                                                                                                                                                                                                                  /                                                                                                                                                                                                                 .                                                                                                                                                                                                       	             1                                                                                                                                                                                            	        -                                                                                                                                                                                                                              0                                                                                                                                                                                                                  0            
                                                                                                                                                                                                                  0                                                                                                                                                                                                                       .                                                                                                                                                                                                                      /                                                                                                                                                                                                                    
 /                                                                                                                                                                                                              -                                                                                                                                                                                                          
       
  .                                                                                                                                                                                                                        0                                                                                                                                                                                                               	    	     -                                                                                                                                                                                                                     .                                                                                                                                                                                                               #               .     	                	           
                                                                                                                                                                                           .                                                                                                                                                                                                                    /                                                                                                                                                                                                                    -                                                                                                                                                                                                                 .                                                                                                                                                                                                                            .                                                                                                                                                                                                             .                                                                                                                                                                                                           /                                                                                                                                                                                                                0                                                                                                                                                                                                             /                                                                                                                                                                                                    	                   0                                                                                                                                                                                                  0                                                                                                                                                                                           	                          /                                                                                                                                                                                                                                        /                                                                                                                                                                                                       
                1                                                                                                                                                                                                          	-                                                                                                                                                                                                             	     	   .                                                                                                                                                                                                                       /                                                                                               
                                                                                                                          0                                                                                                                                                                                           	                            .                                                                                                                                                                                                                           -                                                                                                                                                                                                    .                                                                                                                                                                               
                                      ,          	                                                                                                                                                                                                             0                                                                                                                                                                                                           	    .                                                                                                                                                                                                                  .                                	                                                                                                                                                                                   	                  ,             	                                                                                                                                                                                                                       0                                                                                                                                                                                                              -                                                                                                                                                                                                                                  /                                                                                                                                                                                                                        .          	   
                                                                                                                                                                                              	         2                                                                                                                                                                                                                  -       
                                                                                                                                                                                                      0                                                                                      	                                                                                                                              ,                                                                                                                                                                                                                       -                                                                                                                                                                                                          0                                                                                                                                                                                                                      .                                       '                                                        
                                                                                                                                      /                                                                                      	                                                                                                                                  .                                                                                                                                                                             	                                 0                                                                                                                                                                                                                     -         	                                                                                                                                                                                                                     ,                                                                                   
                                                                                                                         ,                                                                                                                                                                                                            /                                                                                                                                                                                                                       -                                                                                                                                                                                                                                       -                                                                                                                                	                                                                                      .                                                                                                                                                                                                                        -                                                                                                                                                                                                                         -                                                                                           
                                                                                                                      
              /                                    	                                                         	                                                                                                                                    -                                                                                                                                                                                                                     2                                                                                                                                                                                                               /                                                                                                                                                                                                                   1                                                                                                                                                                                         	                           .                                                                                                                                                                                                                       .                                                                                                                                                                                                                             -                                                                                                                                         	                                                                                         ,                                                                                                                                                                                                    .                                                                                                                                   
                                                     
                                 .               	                                                                                                                                                                                                        ,                                                                                                                                                                                                                  	       !                 ,                                                                                                                                                                                                                   /                                                                                                                                                                                                           !             /                	                                                                                                                                                                                                          -                                                                                                                                      
                                                                
                 	  -                                                                                                                                                                                                                             -                                                                                          	                                                                                                                                       .  
                                             	                                                                                                                                                                           .                                                                                                                                                                                                            ,                                                                                                                                                                                                                             0                                                                                                                                                                                                            .                                                                                                                                                                                                                           -                                                                                         	 	                                                                                                                                          .                                                                                                                                                                                                                                 .                                                                                                                                                                                                                 .                                                                                                                                                                                                                             	    ,                                                                                                                                                                                                              	       .        
                                                                                                                                                                                                                 0                                                                                                                                                                                                           
        0                                                                                                                                                                                                                         /                                                                                                                                                                                                             ,                                                                                                                                                                                                                            ,                                                                                  	                                                                                                                           .           	                                                                                                                                                                                                              -                                     5                                                                                                                                                                                                 /                                	                                                      	                                                                                                                                    0                                                                                                                                                                                                        /                                                                                                                                                                                                                    -           	                                                                                                                                                                                	                                    -            
                                                                                                                                                                                                            /                                                                                                                                                                                                                .                                                                                                                                                                                                                 .     	                                                                                                                                                                                                                          	       0                                                                                                                                                                                                                      /                                   	                                                      

                                                                                                                   	              .    
                                                                                                                                                                                                                   /                                                                                                                                                                                                                                .                                                                                                                                                                                                                          /                                                                                                                                                                                                                    1                                                                                                                                                                                                                 /                                                                                                                                                                                        	                           0                                                                                                                                                                                                                        ,                                                                                                                                                                                                                          .                                                                                                                                                                                                                       .                                                                                                                                                                                                                               .                                                                                                                                                                                                              0                                                                                                                                                                                        
                                .                                                                                                                                                                                                                           /                                                                                                                                                                                                                                0                	                                                                                                                                                                                         /                                                                                                                                                                                                                  /                               	                                                                                                                                                                                       -                                                                                                                                                                                                                    
      	       /                                                                                                                                                                                                                            -                                                                                                                                                                                                                           - 
                                                                                                                                                                                                                               -                                                                                                                                                                                         	                          
      .                    	                                                                                                                                                                                                         -                                                                                                                                                                                                         0                                                                                                                                                                                   	                                     0                                                                                                                                                                                                                       -                                                                                                                                                                                                                                          0                                                                                                                                                                                                                 0              	                                                                                                                                                                                                               
   .                                                                                                                                                                                                                  ,           	                                                                                                                                                                                                                     .                                                                                                                                                                                                                 /        
                                                                                                                                                                                                               /                                                                                                                                                                                                                        ,                                                                                                                                                                                                            	               -                                                                                                                                                                                                              0                                                                                                                                                                                                                          ,                                     1                                                        	                                                                                                                                       1                                                                                                                                                                                                                   .                                                                                                                                                                                                            /                                                                                                                                                                                                               -                                                                                                                                                                                                                         
   ,                                                                                                                                                                                                                      -                                                                                                                                                                                                                      -                                                                                                                                                                                                                  .                                                                                                                                                                                                                                 	     .                                                                                                                                                                                                                   0                                                                                                                                                                                                                             .                                                                                                                                                                                                                        -                                                                                                                                                                                                                    0                                                                                                                                                                                                                               -                               
                                                                                                                                                                                     1                                                                                                                                                                                      
                              0                                                                                                                                                                                                             	0                                                                                                                                                                                                                      	  ,                                                                                                                                                                                                                              -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                              
    1                                                                                                                                                                                                           
-                                                                                                                                                                                                                    .              	                                                                                                                                                                                                            -                                                                                                                                                                                                                      	    -           	                                                                                                                                                                                                             -                                                                                                                                                                                                                   -                                                                                                                                                                                                                              -                                                                                                                                                                                                                                
  0                                                                                                                                                                                                                   -                                                                                                                                                                                                                        
  .                                                                                                                                                                                                                              /                                                                                                                                                                                       
                           	           .                                                                                                                                                                                                                         ,                                                                                                                                                                                                             	                         /         /                                                                                                                                                                                                                  .                                    	                                                                                                                                                                       
             .                                                                                                                                                                                                                      -                                                                                                                                                                                                                     	   .                                                                                                                                                                                                                          .                                                                                                                                                                                                              -              	                                                                                                                                                                                                  -                                                                                                                                                                                                        
              	  .                      	                                                                                                                                                                                         	             .                                                                                                                                                                                                                /                                                                                                                                                                                                                     ,                                                                                                                                                                                                                             3             .                                                                                                                                                                                                                      -                                                                                                                                                                                                   -                           	                                                                                                                                                                                  .                
                                                                                                                                                                                                          .                    
                                                                                                                                                                                                      -                                                                                                                                                                                                                      	     .                                                                                                                                                                                                                      .                                                                                                                                                                                                          -                                                                                                                                                                                                                                    -                                                                                                                                                                                                                      
           ,              	                                                                                                                                                                                                       /                                                                                                                                                                                                         /                                                                                                                                                                                                              ,                                                                                                                                                                                                                      .                                                                                         	                                                                                                                       0                                                                                                                                                                                                                        3                                                                                                                                                                                                                  3                                                                                                                                                                             
                              0                                                                                                                                                                             	                                .                                                                                                                                                                                                              2                                                                                                                                                                                                        .                                                                                                                                                                                                                             /                                                                                                                                                                                      
                            .                                                                                                                                                                                                            ,                                                                                                                                                                                                                   /                                                                                                                                                                                                                                    2                                                                                                                                                                                                                       1                                                                                                                                                                                                         /       	                                                                                                                                                                                                                   .                                                                                                                                                                                                                  .                                                                                                                                                                                                               ,                                                                                                                                                                                                                            .                                                                                                                                                                                                                         /                                                                                                                                                                                                                    0                                                                                                                                                                                                                  ,                                                                                                                                                                                                       
                            4       .                                                                                                                                                                                                                     -                                       	                                                                                                                                                                             	               /                                                                                                                                                                                                                          -                                                                                                                                                                                                         	                   
 .                                                                                                                                                                                                                               .                                                                                                                                                                                                                    -                                                                                                                                                                                                                     -                                                                                                                                                                                                            
    	    
  .     	            	                                                                                                                                                                                                             /                                                                                                                                                                                                                   /                                                                                                                                                                                                                      ,                                                                                                                                                                                                                           .                 .                                
                                                                                                                                                                                           .                                                                                                                                                                                                  	       .                               	                                                                                                                                                                               -                                                                                                                                     	                                                                                /                           	                                                                                                                                                                                        .                                                                                                                                                                                                            
               .                                                                                                                                                                                                                  -                                                                                                                                                                                                        .                                                                                                                                                                                                                              .                                                                                                                                                                                                            	                 	   -                                                                                                                                                                                                                 0                                                                                                                                                                                                           .                                                                                                                                                                                                                    -                                                                                                                                                                                                                   /                                                                                           
                                                                                                                  	              .                                                                                                                                                                                                                              0                                                                                                                                                                                                               0                                                                                                                                                                                                       /                                                                                                                                                                                                        -                                                                                                                                                                             	                               /                                                                                                                                                                                                      /                                                                                                                                                                                                                     &        -                                                                                                                                                                                                               ,                                                                                                                             
	                                                         
                                  ,       
     	                                                                                                                                                                                                         /                                                                                                                                                                                                           
      	              0                                                                                                                                                                                                        	              	   0                                                                                                                                                                                                 .        	          	                                                                                                                                                                                                      1                                                                                                                                                                                                           ,              	                                                                         	                                                                                                                            -                                                                                        
                                                                                                                                            -  	                                                                                                                                                                                                                         ,                                                                                                                                                                                                    ;                                      .                                                                                                                                                                                                                      .                                                                                                                                                                                                                            
  /                 	                                                                                                                                                                                                               -                                                                                                                                                                                                                                 -             	                                                                                                                                                                                                               ,                                                                                                
                                                                                                                   
                       -              
                                                                                                                                                                                                       /                                                                                                                                                                                                                   -              	                                                                                                                                                                                                               ,                                                                                                                                                                                                                                1                                                                                                                                                                                                                                  .                                                                                                                                                                                                               
                   -                                                                                                                                                                                                                     -                                                                                                                                                                                                             
              
 -                             
                                                                                                                                                                                                .                                                                                                                                                                                                                    -                             	                                                                                                                                                                                                    -                                   	                                                                                                                                                                	           -          
                                                                                                                                                                                                               .                                                                                                                                                                                                                          .                                                                                                                                                                                                                  0                                                                                                                                                                                                                      -                                                                                                                                                                                                                             ,        
                                                                                                                                                                                                                                    -      	     
                                                                                                                                                                                                                       .                                                                                                                                                                                                                    .                                                                                                                                                                                                      -                                                                                                                                                                                                                         .                                                                                                                                                                                                                            .                              
                                                                                                                                                                                             .                                 	                                                                                                                                                                                            .                                                                                                                                                                                        	                         /                                                                                                                        	                                                                                   .                                                                                                                                                                                                                  .                                                                                                                                                                                                              -                                                                                                                                                                                                	                                        /                                                                                                                                                                                                             	.                                                                                                                                                                                                                     .                                                                                                                                                                                                                 .                                                                                                                                                                                                          
                    
     /                                                                                                                                                                                                                   /              
       	                                                                                                                                                                                                            /                                
                                                                                                                                                                                   -                                                                                                                                                                                                                          	  -                                                                                                                                                                                                                  -                                                                                                                                                                                                                    -                                                                                                                                                                                                                             .                                                                                                                                                                                                                                      .        
                                                                                                                                                                                                              -                                                                                                                                                                                                              	                   0                                                                                                                     
                                                                                        .                                                                                                                                                                                                                      -                                                                                                                                                                                                                             ,                                                                                                                                                                                                                               $	             .                                                                                                                                                                                                                             .                                                                                                                                                                                     	                              /               

                                                                                                                                                                                          	                 -                                                                                                                                                                                                                                           ,                                                                                                                                                                                                                               	     0                                                                                        	                                                                                                                             0                                                                                                                                                                                                                -                                                                                                                                                                                                                              /      	                            
                                                                                                                                                                                .                                                                                                                                                                                                                   -                                                                                                                                                                                                                         /                                                                                                                                                                                                               -                            	                                                                                                                                                                                               .                                                                                                                                                                                                                            
    -                                                                                                                                                                                                                          .                                                                                                                                                                                                                      - 
                                                                                                                                                                                                                       -                                                                                                                                                                                                                                ,                       	                                                                                                                  
                                                                                            .                                                                                                                                                                                                        
           0                                                                                                                                                                                                            -                                                                                                                                                                                                                                    	.                                                                                                                                                                                                                                    .                                                                                     
                                                                                                                                  1                                                                                                                                                                                                                    0                                                                                                                                                                                         
                            /                                                                                                                           	                                                                                    .                                                                                                                                                                                                                   .                                                                                                                                                                                 
                               -                 	                                                                                                                                                                                                                 /                                                                                                                                                                                                     .                                                                                                                                                                                                          	           -                                                                                                                         
                                                                                              -                                                                                                                                                                                                             	                     	    .                                                                                                                                                                                                                     .    	                  	                                                                                                                                                                                                         .      	                                                                                                                                                                                                                  ,                                                                                                                                                                                                                    "             -                                                                                                                                                                                                           -                                                                                          	                                                                                                                                         -                   	                                                                                                                                                                                                      -                                                                                                                                                                                           +                            
       -                                                                                                                                                                                                                      .                                                                                                                                                                                                                     .           	                                                                                                                   	                                                                                             -                                                                                                                                                                                                                        -                                                                                                                                                                                                            	                 ,                                                                                                                                                                                                                              (
              .                                                                                                                                                                                                                             .                                                                                                                                                                                                                     -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                    
                     -                                                                                                                                                                                                                                   /                                                                                                                            
                                                                           
                  /      	                                                                                                                                                                                                      /                                                                                                                                                                                                                               /      	                                                                                                                                                                                                                .                                    
                                                                                                                                                                                -                                                                                                                                                                                                                        .                                                                                                                                                                                                          .                                                                                                                                                                                                                         /                                                                                                                                                                                                                           	  /                                                                                                                                                                                                                              .                                                                                                                                                                                                                           .     	               	                                                                                                                                                                                                         -                                                                                                                                                                                                                                  ,                      
                                                                                                                  	                                                                                                  -                                                                                                                                                                                                               
      .                                                                                                                                                                                                        /                                                                                           	                                                                                                                          0                                                                                                                                                                                                                	             /                                                                                                                                                                                                                                .                                   	                                                    
 
                                                                                                                                 /                                                                                                                                                                                            
                         .                                                                                                                                                                                                          -                                                                                                                                                                                                                -                                                                                                                                                                                                           .                                                                                                                                                                                                                          )         ,                                                                                                                                                                                                                   .                                                                                                                                                                                      	                              .             	                                                                                                            
                                                                                           ,                                                                                                                                                                                                         
          	         /                               	                                                                                                                                                                                     -                                                                                                                                                                                                                  %                  /   
                                                                                                                                                                                                                   /                                                                                                                                                                                                                                  .                                                                                                                                                                                                           .                                                                                      	                                                                                                                             -    	                                                                                                                                                                                                                         .                                                                                                                                                                                                         	                               -                                                                                                                                                                                                                                    ,                                                                                                                                                                                                               ,                                                                                                                                                                                                     	                            %          ,                                                                                                                                                                                                                                  -              	                                                                                                                                                                                                             -                                                                                                                                                                                                                            /                                                                                                                                                                                                                             (          -                                                                                                                                                                                                                               	  .                                                                                                                                                                                                                      .                      	              	                                                                                                                                                                                      .                                                                                                                                                                                                                                 -                                                                                                                                                                                                                             7                 ,                                                                                                                                                                                                                                        .                                                                                                                                                                                                        ,                                                                                                                                                                                                                   !            
    ,                                                                                                                                          
                                                                                     
      -                                                                                                                                                                                                                                             -                                                                                                                                                                                                   	                                    -                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                     
 -                                                                                                                                                                                                                                     .                                                                                                                                                                                                                                  .                     
                                                                                                                                                                                                         ,                                                                                                                                                                                                                                   -                                                                                                                                                                                                                             /                                	                                                                                                                                                                                   0                                                                                                                                                                                                                        ,                                                                                                                                                                                                     	    
                           ,                                                                                             	                                                                                                                                   .                                                                                                                                                                                                                                  -                                                                                                                                                                                                                  ,                                                                                             
                                                                                                                               ,                                                                                                                                                                                                                                   0                                                                                                                              
                                                      
                              /                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                  .          $                                                                                                                                                                                                                   .                                                                                                                                                                                                                        	          
   ,                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                  ,               	                                                                                                                                                                                                                   -                                                                                                                                                                                                                                /                                                                                                                                                                                                                                -               )                                                                                                                                                                                                                   ,                   	                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                                --                                                                                                                                                                                                                     
    	          -                                                                                                                                                                                                                               ,                                    
                                                                                                                                                                                    ,                                                                                                                                                                                                                               !       -                                                                                                                                                                                                                           -                                                                                                                                                                                                                          -           ,                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                    !     .                                                                                                                                                                                                                     
    ,                                                                                                                                                                                                                                                     -                      	                                                                                                                                                                                                              ,                 
                                                                                                                                                                                                               -                 	                                                                                                                                                                                                               
      -                                                                                                                                                                                                                              .                                	                                                         
                                                                                                                                      /                                                                                                                                                                                                                       -                                                                                                                                                                                                                     	      -                                                                                                                                                                                                                      -               
                                                                                                             	                                                                                            ,                                                                                                                                                                                                                          -        
                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                              ,                    0                                                                                                                                                                                                                       -                                                                                                                                                                                                                                      -                
                                                                                                                                                                                                            ,                                                                                                                                                                                                                                 &              ,            	      (                                                                                                                      	                                                                                                       ,                                                                                                                                                                                                                                         -         %                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                      	            ,                                                                                             !                                                                                                                                         ,                                   )                                                                                                                                                                                                             ,                                       #                                                                                                                                                                                                ,                                                                                                                                                                                                          	                                     ,                                                                                                                                   #                                                                                        -                                                                                                                                         -                                                                                                ,                                                                                                                                           )                                                                                                   ,                                                                                                                                                                                                                                     (           ,            (                           	                                                                                                                                                                                                         ,                                                                                                                                                                                                                          	              .               
                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                           ,          !                                                                                                                                                                                                                          -                                                                                                                                                                                                              %               /         	             
                                                                                                                                                                                                         ,                                                                                                                                                                                                                                      -                                                                                                                                                                                                                           
.                                                                                                                                                                                                            
              -                                                                                                                                                                                                                                   .                                                                                                                                                                                                                               	      ,                 		                                                                                                                                                                                                                .                                                                                                                                                                                                                -                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                            -                                                                                                                                                                                                                  
      
        ,                       
                                                                                                                                                                                                       .                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                   
            	  -                   	                                                                                                                                                                                        	                        ,                                                                                                                                                                                                                                                /                                                                                                                                                                                                                                              /                                                                                                                                                                                                                                ,                                                                                       	                                                                                                                                        -                                                                                                                                                                                                              ,                                                                                                                                                                                                                                 
     ,                                      $                                                                                                                                                                                                  .                                                                                                                                                                                                                                .                                                                                                                                                                                                                      ,                                	                                                                                                                                                                                                ,                                                                                                                                                                                                                                     $         ,                                                                                                                                                                                                                                           ,                                                                                                                                                                                                         	                       $   	     /                      
                                                                                                                                                                                                       -                                                                                                   	                                                                                                                         
                  ,                                                                                                                                                                                                                                        ,                                                                                                                                                
                                                         
                	           
      -      	             	           	                                                                                                                                                                                                  ,                                                                                                                                                                                                                                           
      ,                                       
                                                                                                                                                                                                  ,                                                                                                                                                                                                                                  /                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                                   .                                                                                                                                                                                                                          .                                                                                                                                      '                                                                                               ,                                                                                                                                                                                                                                              -               	                                                                                                                   	                                                                                          -                                                                                                                                        
                                                                                   -                                                                                                                                     	                                                                                       -                                                                                                                                                                                                              !             
     -                                                                                                                                                                                                                    -                                                                                                                                                                                                                          	   ,                                                                                                                                                                                                                                  	   ,                                                                                                                                         	                                                                                          -                                                                                 
                                                                                                                                 ,                                                                                                                                                                                                                    	            .                                                                                                                                                                                                                          -                                                                                                                                                                                                                          	  -                                  	                                                                                                                                                                                      ,                                                                                                                                                                                                                     -                                                                                                                                                                                                      	                          '      ,                                                                                                    
                                                                                                                                    -                                                                                                                                                                                                            	              ,                         	                                                                                                                                                                                                            -                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                           -                               	                                                                                                                                                                                               -                                                                                        	                                                                                                                                      -                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                     -                                                                                                                             	                                                                                                 .              	                 	                                                       
                                                                                                                                      -                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                      -                                                                                                                                                                                                                          	             ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                             
       &          ,                                                                                                                                                                                                                                          -                                                                                                                                                                                                                   
         	   ,                                                                                                                                                                                                                       
                 ,                                                                                                                                                                                                                          8                     ,                 $                                                                                                                                                                                                                           .                                                                                                                                                                                                                   
               -       	                          	                                                                                                                                                                                          -                                                                                                      	                                                                                                                                  -                                                                                           
                                                                                                                               /                                                                                                                                                                                                                         0                                  -                                                                                                                                                                                           ,                                                                                                                                                                                            	                                 ,                                                                                                                                                                                                               
                ,                                                                                                                                                                                                                              ,                                         '                                                                                                                                                                                                        ,                                                                                                                                                                                                                                    #               ,                     	                                                                                                                                                                                                	       ,                                                                                                                                                                                                                                     -                
                                                                                                               	                                                                                           -                                                                                                                                                                                                                                                ,                                        
                                                                                                                                                                                                     -                                                                                                                                                                                                                	                  ,                #                                                                                                                                                                                                                      ,                                                                                                                                                                                                                     
             ,                                                                                           	 	                                                                                                                                                  ,                                      	                                                                                                                                                                                  "                    ,                       
                                                                                                                                                                                              
                     ,                                                                                                                                                                                                 &                                   -                                 
                                                                                                                                                                                      
      -                                                                                                                                                                                                                        ,                                                                                                                                                                                                                              )           ,                                                                                                                                                                                                                                 	       ,              	                                                                                                                                                                                                            	            ,            	                                                                                                                            	                                                                                            -                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                '     
    -                                                                                                                                                                                                                               
             ,                                       	                                                                                                                                                                                                   -                 
                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                     ,                                                                                             %                                                                                                                          	                 -                                                                                                                                                                                                                           .                                                                                                                                                                                                                      (             ,                                                                                                                                                                                                                       ,                                      !                                                                                                                                                                                       ,                                     D                                                                                                                                                                                                           ,                                     +                                                                                                                                                                                                              ,                                     0                                                        	                                                                                                                                            ,                                                                                                                                                                                                                                                 ,            	                                                                                                                                                                                                                    -                                                                                                                                                                                                                                 ,                                          "                                                                                                                                                                                             
            -                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                      	      -            ,            
                                                                                                                                                                                                                 ,                                      
                                                                                                                                                                                            ,               	                                                                             %                                                                                                                                                  -                                                                                                                                                                                                                                          -                            $                                                                                                                                                                                                     ,                                                                                                                                                                                                    	 
                               ,                                                                                                                                                                                                           '                                     .                                                                                                                                                                                                                                     ,                                                                                                                                                  G                                                                                                     ,                                                                                                                                                                                                                                      	   	         ,                                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                              &       ,                                                                                                                                                                                                                                   -                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                               ,                                                                                                                                                                                                                               -               =                                                                                                                                                                                                                           -                                                                                                                                                                                                                            -                                     
                                                                                                                                                                                       ,                                     	                                                                                                   
                                                                                                      ,                                                                                                                                                                                                                                     -                                                                                                                                                                                                                            	       ,                  
                                                                                                                                                                                                                  -                                                                                                                                                                                                                    -                                                                                                                                                                                                                        
     $              ,                                                                                                                                                                                                                                                  -                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                          	,            
                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                            -                                                                                                                                                                                                                                    ,               
                                                                                                                                                                                                           ,                                                                                                                                                                                                                                              -                                                                                                  +                                                                                                                                      ,                                                                                                                                                                                                                                   ,                 
                                                                                                                                                                                                            .                                                                                                                                                                                                                             %                   -                                    &                                                                                                                                                                                                         ,                                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                      ,             	                                                                                                                                                                                                                             ,                                      
                                                                                                                                                                                             ,             1              
                                                                                                                                                                                                                -                                                                                                                                                                                                                          -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                     ,                                                                                                                                          
                                                                                             -                                 	                                                                                                                                                                                       ,             <                           
                                                                                                                                                                                                          ,                                                                                                                                                                                                                                     ,                         	                                                                                                                                                                                                               ,                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                     -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                            ,                   	                                                                                                                         -                                                                                                -                	                                                                                                                                                                                                                ,                                                                                                                                                                                                                                              .                                                                                               	                                                                                                                                    -                                                                                                                                                                                                                                         ,                                                                                           	                                                                                                                                    ,                                                                                                                                                                                                                                                     .                                                                                                                                                                                                                              -                                                                                                                                                                                                                                  ,      	                 
                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                       -                                                                                                                                                                                                                           	      2           -                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                      !                 ,                                                                                                                                                                                                                                     .                                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                           -                                                                                                                                                                                                                                            ,                                                                                             
                                                                                                                                  .                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                           
 ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                               	                                  ,       
                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                             ,                          
                                                                                                                           	                                                                                            /                                                                                                                                                                                                                     ,                 %                                                                                                                                                                                                                                /                                                                                                                                                                                                                                  -                   *                                                                                                                                                                                                                       ,                                                   	                                                                                                                                                                               ,                                 	                                                           	 
                                                                                                                                              ,                                                                                                                                                                                                                         -                      
                                                                                                                                                                                                        ,               
       
                                                                                                                                                                                                               ,                                                                                                                                                                                                                                     -                                                                                                                                                                                                                                         ,                                 +                                                                                                                                                                                                   ,                                                                                                                                                                                                                                         -                                                                                                                                       	                                                                                                 ,                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                                    
-                                                                                                                                                                                                                                       ,                        	                                                                                                                                                                              	                                       -                                                                                                                                                                                                                                        ,                                                                                                                                             #	                                                                                                   ,              	       
                                                                                                                                                                                                  -          %                                                                                                                                                                                                                                /                                                                                                                                                                                                                    #              ,            &              
                                                                                                                                                                                                                        -                                                                                                                                                                                                                                 ,                '                                                                                                                                                                                                                          -                                                                                                                                                                                                                             "            ,            .                                                                                                                                                                                                                                          ,                                                                                                                                                                                                       )                            	      ,                                                                                                                                        	                                                                                      ,                                                                                                                                                                                                                    
             .                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                         	                -             
       	                                                                                                                                                                                                                 ,                                                                                           	                                                                                                                               -                                                                                                                                                                                                                     &                ,                                                                                                                                                                                                                                  -                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                      -                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                    ,                 
                                                                                                                                                                                                                 
     .                                                                                                                                                                                                                         -                                                                                                                                                                                                                               -                	                                                                                                                                                                                                                      -         #                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                           (           	   ,                  (      
                                                                                                                                                                                                   	                 -                                                                                                                                                                                                                                      -                                                                                                                                                                                                                          	     -                                                                                                                                                                                                                              2           	     ,                                                                                                                                                                                                                                       -                                                                                                                                                                                                                ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                  
              ,                                                                                                 4                                                                                                                            	               ,          
                                                                                                                                                                                  
                                      /                                     1                                                                                                                                                                                                          ,                                                                                                                                                                                                            
                 
                -                                                                                                                                                                                                                                 -                                                                                                                                                                                                                           /                                                                                                                                   )                                                                                                    ,                                                                                                                                                                                                                                           ,                      
                                                                                                                                                                                                             -                                                                                                                                                                                                                           -                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                 "            -                                                                                                                                                                                                                                              .                                                                                                                                                                                                                      	             ,                                                                                                                                                                                                                                     -                                                                                                                                                                                                                   !              ,           
                          
                                                                                                                                                                                 	                  .                                                                                                                                                                                                                       #              -     	                                                                                                                                                                                                                          -                                                                                                                                           	                                                                                             ,                                                                                                                                       
                                                                                         -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                             ,                                       
                                                                                                                                                                                          -                    
                                                                                                                                                                                                              ,                                                                                                                                                                                                                                    
      ,                                                                                                                                                                                                                  	          ,                                                                                                 
                                                                                                                          (                   -                                                                                                                                                                                                                        ,                                                                                                                                                                                                                      .                       	                                                                                                                                                                                                             -                                                                                                                                                                                                 
                 
            ,                      
                                                                                                                                                                                                           /                                                                                                                                                                                                                        -                                                                                         
                                                                                                                                     ,                                     	                                                                                                                                                                                                     ,                    	                                                                                                                                                                                                        .                                                                                                                                                                                                                               +   	      ,                                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                       ,                 
                                                                                                                                                                                                                         -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                      	-                                        	                                                                                                                                                                                        -                                                                                                                                                                                                                             
            /                                                                                                                                 	                                                                                        ,                                                                                                                                                                                                                          ,                                                                                            	                                                                                                                                    	.                                                                                                                                                                                                                      
            ,             	                                                                                                                                                                                                                          -                                 	                                                                                                                                                                                                        ,                        
                                                                                                                                                                                                                   -                                                                                                                                                                                                                                        /                                                                                                                                                                                                                      -                                   	                                                                                                                                                                                        ,    	                                                                                                                                                                                                                                           .                                                                                                                                                                                                                             -        
                      	                                                                                                                                                                                           -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                               .                                                                                         
                                                                                                                                       .             
                                                                                                                                                                                                       -                                                                                                                                                                                                                       -                                                                                                                                                                                                                              -                                                                                                                                                                                                                 	                 .                                                                                            	                                                                                                                                 -                                                                                                                                                                                                #                                  ,                                   	                                                                                                                                                                                              -                                                                                                                                                                                                                   -                                                                                                                                                                                           
                                	    ,                                                                                                                                                                                                                                          0                                                                                                                                                                                                                          -               
                                                                                                                                                                                 
                            -              
                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                 -                      
                                                                                                                                                                                                                 -                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                      -                                                                                                                                                                                                                         -                                                                                                                                                                                                                             -                                                                                                                                                                                                                            -                                                                                             	                                                                                                                           	                 ,                                                                                                                                                                                                                         ,                                                                                                                                                                                                              ,                                                                                                                                                                                     
                                 .                                                                                                                              
                                                                                                -      	                                                                                                                                                                                                                           /                                 
                                                                                                                                                                                                 .                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                     ,                                      	                                                                                                                                                                                              .                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                 -            ,           '                                                                                                                                                                                                                        ,          
             
                                                                                                                                                                                                           ,                                                                                                                                                                                                                                        ,                                                                                      	                                      	                                                                                          .                                                                                                                                                                                                                            ,          	                                                                                    
                                                                                                                                      	,                                                                                                                                                                                                   	                                .                                                                                                                                                                                                                      -                                                                                                                                                                                                 
                                  ,                                                                                                                                                                                                                               	   /                                                                                                                                                                                                                       	         -                                         	                                                           
                                                                                                                                 ,                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                 .         &                                                                                                                                                                                                                    	         ,                                                                                                                                                                                                                                            .                      
                                                                                                                                                                                              	              ,                                                                                                                                    
                                                                                                     -                                                                                                                                                                                                                        ,                                                                                                
                                                                                                    	                           -                                                                                                                                                                                                                                         .                                	                                                                                                                                                                                       -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                       .                                                                                                                                                                                                                      ,                                                                                                     
                                                                                                                                        -                                                                                                                                                                                                                                          -                                                                                                  	                                                                                                             
              ,                                                                                                                                                                                                                             ,                  
                                                                                                                                                                                                            .                    	                                                                                                                                                                                                                       -                                                                                                                                                                                                                          -                                                                                                                                                                                                                      
     
          ,                                                                                                                                                                                                                 	                   ,                                                                                           	                                                                                                                                       .                                                                                                                                                                                                                      .             	                                                                                                                                                                                                                   -                                                                                                                                                                                                                         
.                                                                                                                                                                                                                            0                            	                                                                                                                                                   	                                 .                                                                                                                                                                                                                             /                                                                                                                                                                                                       -      	     "                                                                                                                                                                                                                                -                                                                                                                                                                                                                      -          
                                                                                                                                                                                                         ,                                   %                                                                                                                                                                                                      ,                                                                                                                                                                                                                                      0                                                                                                                                                                                                                                -                                                                                                                                                                                                                         ,                          	              	                                                                                                                                                                                                 -           
                                                                                                                                                                                                                           ,                                                                                                                                                                                                                   -                             
                                                                                                                                                                                     ,                                                                                                                                                                                                                         -                                                                                                                                                                                                                                     -                                                                                                                                                                                                                     .                                                                                                                                                                                                               ,                                                                                                                                                                                                             
   	         -                                                                                                                                                                                                                                 .                                                                                                                                                                                                                                ,                                                                                                                                                                                                                          ,                                                                                                                                           

                                                                                   	   .                   
                                                                                                                                                                                                              /                                                                                                                                                                                                                    ,                      
                                                                                                                                                                                                               -                                                                                                                                                                                                                          -                                                                                                                                                                                                                           .                                                                                                                                                                                                    
               -                                                                                                                                                                                                            -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                  
-                                                                                                                                                                                                                       	  .                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                             	       -                	                                                                                                                                                                                                                 ,            	                                                                                                                               	                                                                                           -      
                                                                                                                                                                                                                                	             ,                                                                                                                                                                                                                                      -          	                                                                                                                                                                                                                   .                                                                                                                                                                                                                 -                                                                                                                                                                                                                         	                 -                                                                                                                                   
                                                                                    ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                
-                                                                                                                                                                                                                                   	              -                                                                                                                                                                                                                                        .                            	                                                                                                                                                                                            ,                                                                                                                                                                                                                              ,                )                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                    >	                    .                      
                                                                                                                                                                                                                -                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                    ,                                                                                                      
                                                                                                                                             ,                             
                                                                                                                                                                                       -                                                                                                                                                                                           
                         -                                                                                                                                                                                                                        ,                                                                                                                                                                                                           	                           	    -                                                                                                                                                                                                                          -                                                                                            
                                                                                                                                   0                                    4                                                                                                                                                                                                   ,                                                                                                                                                                                                                           
            -                                                                                                                                                                                                                   
      -                                                                                                                                                                                                                         -                                                                                                                                        ;                                                          	                                      ,                                                                                                                                                                                                                                           3          -                                                                                                                                                                                                          	       .                                                                                                                                                                                                	                       
           ,                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                   
       0          ,       -                         
                                                                                                                                                                                                         .                                                                                                                                                                                                                 	               ,           #            
                                                                                                                                                                                                                       -                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                  -                                                                                                                                                                                                                     !              ,                        	                                                                                                                                                                                                       ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                   
-                                                                                                                                                                                                                       	                    ,         
   	       
                                                                                                                                                                                                                 /                                                                                                                                                                                                                                         ,            	             	                                                                                                                            	                                                                                   -                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                                       .                                                                                                                                                                                                                                  7             ,                                                                                                                                                                                                                                          -                        	                                                                                                                                                                                                              
       -                                                                                                                                                                                                                         -                                                                                                                                                                                                                                  ,            	                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                     -               	                                                                                                                                                                                                                      -                                                                                                                                                                                                            	                 .                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                           9      	      .                #                                                                                                                                                                                                                          -                                                                                                                                                                                                                                     G              ,            	           	                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                               ,              )      	                                                                                                                                                                                                                      -                                                                                                                                                                                                                                    	     ,           (     	                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                    2                   ,                                                                                                                                                                                                                                            ,                                     $                                                                                                                                                                                                  -                                     	                                                                                                                                                                                             ,                                                                                                      	                                                                                                      (                                 ,                                                                                                                                                                                                              +                           
      ,                                                                                                                                            	                                                                                   	          -                                                                                                                                                                                                                        ,                                                                                                                                                                                                                
                                  ,                  

                                                                                                                                                                                                                          -                                                                                                                                                                                                                 0                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                           <          -           /     	                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                            -                       	                                                                                                                                                                                          
              ,                                                                                                                                                                                                                          
             "            ,                 /                                                                                                                          	                                                                                                    /                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                            -                                                                                               
                                                                                                                          	  -                                 
                                                           
                                       	                                                                                          .                                                                                                                                                                                                                              .                                                                                                                                                                                                                                ,                                                                                                                                                                                                                             ,                                                                                                                                                                                                                       	    .                                                                                                                                      	                                                                                             .                                                                                                                                                                                                                                    -                                                                                          	                                                                                                                          ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                            .          
                                                                                                                                                                                                                    -                                                                                                                                                                                                                               .                                                                                                                                                                                                                              ,                                                                                                                                                                                                        
                -                                                                                                                                                                                                                             	    ,                                                                                                                                                                                                                            -                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                              
,                                                                                                                                    	                                                                                               -                                                                                                                                                                                                                          .                                                                                                                                                                                              
                                 0          
                                                                                                                                                                                                                          ,                                                                                                                                                                                                                               	  	-                                                                                                                                                                                                                                  -           &                                                                                                                                                                                                                               -                                                                                                                                                                                                                        -                                                                                                                               
                                                                                                ,                                                                                                                                                                                                                              ,                                    	                                                       
                                                                                                                                    ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                	-                                                                                                                                                                                                                                  .                                                                                                                                                                                                                              -                                                                                                                                                                                                                             -                                                                                                                                                                                                                              
-                 
                                                                                                                                                                                                        ,                                                                                                                                    
                                                                                                  ,                                                                                                                                    
                                                        	                              .                                                                                                                                                                                                                                    -                                                                                                                                                                                                             
           -                                                                                                                                                                                                                                1                      
                                                                                                                                                                                                       	     -                                                                                                                                                                                                                      	                ,         	                                                                                                                                                                                                                           -                               	                                                                                                                                                                                             -                                                                                                                                                                                                                                ,                                      
                                                                                                                                                                                               -                                                                                                                                                                                                    (                                  ,                                                                                                                                   	                                                                                                ,                                                                                                                                                                                                                                  -                                                                                                                                                                                                                           -                                 
                                                   

                                                                                                                                   -                                                                                                                                                                                                                             
     -                             	               	                                                                                                                                                                       -                                                                                                                                                                                                                                     
      -                                                                                                                                                                                                
                              -                                                                                                                                                                                                                                              .                                                                                                                                                                                                                     -                                                                                                                                                                                                                                      /                                                                                                                                        
                                                                          
                   ,                                                                                                                                                                                             
                                   .                                                                                                                                                                                                       
                -                                                                                                                                                                                                                                 -                                                                                                                                                                                                                           
      .               
                                                                                                                                                                                                         -                                                                                                                                                                                                                          -                                                                                                                                                                                                                                     .                                                                                                                                                                                                                                      -                 
                                                                                                                                                                                                                     .                                                                                                                                                                                                               -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                             	        ,       	                                                                                                                                                                                                                              /                                                                                       
                                                                                                                               -       	                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                          .                                                                                                                                                                                                                                  ,                                     (   
                                                                                                                                                                                                          ,                      	                                                                                                                                                     
                                                            ,                                                                                                                                                                                                                                          -                                                                                                                                            
                                                          	                             ,                                                                                                                                                                                                                                                   ,                                	                                                                                                                                                                                                      -                                                                                                                                                                                                                                             ,                 
                      
                                                                                                                                                                                                 ,                                       	                                                                                                                                                                      
          
    ,                                                                                                                                                                                                                               .                                                                                                                                                                                                                                      ,           "                                                                                                                                                                                                                           -                                                                                                                                                                                                                         -                                                                                                                                                                                                                              0                                                                                                                                                                                                                         -                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                        .       
                                                                                                                                                                                                                          -                                                                                                                                                                                                                                   ,          	     	              
                                                                                                                                                                                                 -                                                                                                                                                                                                                              .         	                                                                                                                                                                                                          
        -          	                                                                                                                                                                                                     /                                                                                                                                                                                                                                ,         	                                                                                                                                                                                                              0                                                                                                                                                                                                                 
         ,                                                                                                                                                                                                                 .                                                                                                                                                                                                                              #         ,                                                                                                                                                                                                                           .                                                                                                                                                                                                                              	,                                                                                                                                                                                                                                       -                                                                                                                                                                                                                                 -                                                                                                                                                                                                                	-                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                .              
                                                                                                                                                                              
                                    .                                                                                                                                                                                              
                          -                                                                                                                                                                                                   	                                     ,                                                                                                                                                                                               	          	                   
     ,                	                                                                                                                                                                                                                              ,                                                                                                                                                                                                                       	 	   -                  
                                                                                                                                                                                                        .                                                                                                                                                                                                                                   .           
                                                                                                                                                                                                                   /                                                                                                                                                                                                                    .                                                                                                                                                                                                                             -                                                                                        	                                                                                                                                 	,                                                                                                                                                                                                                                 	-                                                                                                                                                                                                                                  -                                     
                                                                                                                                                                                          -                                                                                                                                                                                                   	                            
-                                                                                                                                                                                                    	                            
     	,                                                                                                                                                                                                                                      -                                                                                                                                                                                                                            ,                                                                                                                                                                                                                             
     ,                                                                                                                                                                                                                                     -                                                                                                                                                                                       	                             	     ,           
                                                                                                                                                                                                                 -                                                                                                                                                                                                                      #                ,                 
                                                                                                                  	                                                                                                    -                                                                                                  
                                                                                                                            	     .                                                                                                                                                                                                                         ,                                                                                                                                                                                                                              -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                           .                                                                                                                                                                                                                             -                                   
                                                                                                                                                         
                                    ,                                                                                                                                                                                                                    	.                                                                                                                                                                                                            -                                                                                                                                                                                                                                    ,                                	                                                                                                                                                                                      
,                                                                                                                                                                                                                        
     	,                 
                                                                                                                                                                                                            
/                                                                                                                                                                                                                       	        ,                                                                                                      	                                        	                                                           
                        -         	                                                                                                                                                                                                                              ,                                                                                                                                                                                                                         .                        	                                                                                                                                                                                                           .                                                                                                                                                                                                                                     -                                 
                                                                                                 	                                                                                     .                                                                                                                                                                                                                      .                                                                                                                                                                                                                                   .                                                                                                                                                                                                               ,              	                                                                                                                                                                             	                        
     .                      
                                                                                                                                                                                                                   -                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                       .                                                                                                                                                                                                                   -           	                                                                                                                                                                                                                        -                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                      -                                                                                                                                                                                                                                          /                                                                                                                                                                                                                        	-                                                                                                                                                                                                                                ,                                         
                                                           	                                                                                                                                  ,                                                                                                                                                                                                 	                                .                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                            
      .                                                                                                 	                                                                                                                      
                -                                                                                                                                                                                           	                            ,                                                                                                                                  "                                                                                                 -                                                                                                                                                                                                                                       -                                                                                                                                                                                                                             	   
   .                                                                                                                                                                                                                               ,                     	                                                                     
                                                                                                                                          -                                                                                                                                                                                                                                             /                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                    -                                                                                                                                                                                                                                  .                                                                                                                                                                                                                 .                                                                                                                                                                                                                    ,                                                                                                                                                                                                                       &
             ,                                                                                                                                                                                                                                  .                                                                                                                                                                                                                                        .                                                                                                                                                                                                                                   ,                               
                                                                                                                                                                                         -          	                                                                                                                                                                                                                   -       	                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                     ,                	                                                                                                                   
                                                                                         -                                                                                                                                                                                                                              -                                                                                                                                                                                                                       -                                                                                                                                                                                                                                 "           ,                                                                                                                                                                                                                                      -                      	                                                                                                                                                                                                                  -                                                                                                                                                                                                                                   ,                                                                                                                                                                                                              	            	      /                                                                                                                                                                                                            /                                                                                                                                                                                                                     ,                                                                                                                                                                                                              
       ,                                                                                                                                                                                                                                       ,                                                                                                                                                                                                     	                                -                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                           -               	$                                                                                                                          
                                                                                                  -                                                                                                                                                                                                                               ,                                                                                                                                        	                                                                             
        ,                                                                                                                                                                                                                         	      "            -                                                                                                                                                                                                                                           .         
                                                                                                                                                                                                        
                 -                                    
                                                                                                                                                                                            ,                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                               	         
    ,                                                                                                                                                                                                                                    ,                 	                                                                                                                           "                                                                                                     -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                        	            ,                                                                                                                                                                                                                                     .                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                          -                                                                                                                                                                                                                                                  ,          %   	                	                                                                                                                                                                                                           -                                                                                                                                                                                                                          -                                                                                                                                                                                                               
              ,                                                                                                                                                                                                                               ,       	                                                                                                                                                                                                                             -                                                                                                                                                                                                                    !                ,                                                                                                                                                                                                                                   -                                                                                                                                                                                                           <                                      -                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                        -                                                                                                                                                                                                                                   -                                                                                                                                                                                                                                        -                                                                                                                                                                                                                          
       -                                                                                                                                                                                                                               ,                                                                                                                                                                                                          	                     ,                                                                                                                                                                                                                             -                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                  -                                                                                                                                                                                                                  	               /                                                                                                                                                                                                                                       ,       
                         	                                                                                                                                                                                                    ,                                                                                                                                                                                                                         
.          	     	                                                                                                                                                                                                                     ,                               
                                                                                                                                                                                             ,                                   
                                                                                                                                                                                                   0                                                                                                                                                                                                                        /                                                                                             	                                                                                                                                       .                  	                                                                                                                                                                                                              ,                                                                                                                                                                                                                                   /                                                                                                                                                                                                                        .                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                     -          
                                                                                                                                                                                                                            -                                                                                                                                                                                                           
            /                                                                                                                                                                                                                     ,                                                                                        	                                                                                                                                  ,                                                                                             & 	                                                                                                                                              .                                                                                                                                                                                                                  .                                                                                                                                                                                                                         ,                 	                                                                                                                                                                                                           ,                                                                                                                                                                                                           ' 
                                 .                              	                                                                                                                                                                               
          .                                  	                                                                                               !                                                                                                ,                                                                                                                                                                                                                            0                                                                                                                                                                                                                       .                                                                                                                                                                                                           -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                        .         
                        	                                                                                                                                                                                       	              -                                                                                                                                                                                                                             -                                                                                                                                                                                                                                         ,                                                                                                                                        	                                                                                   .         	                                                                                                                                                                                                                          ,                                                                                                                                                                                                                               .                                                                                                                                                                                                                                ,                                                                                                                                                                                                                              ,           	                                                                                                                                                                                                         	          /                                   	                                                                                                                                                                                  .               	                                                                                                                                                                                                                 ,                                                                                                                                                                                                                       -                                                                                                                                                                                                                               -                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                 -                                                                                                                                                                                                            	          .                                                                                                                                                                                                                                           .                                                                                   
                                                                                                                            ,                                                                                                                                                                                                                                         .                                                                                                                                                                                                         	               -                                                                                                                                                                                                                                   -                                                                                    	                                                                                                                              /                                                                                                                                                                                                                                  .                                                                                                                                                                                       	                          	    -                                                                                                                                                                                                                                 -                                                                                                                                                                                                                             ,                                                                                                                                                                                                      	                                     ,                                                                                                                                                                                                                                     !          ,      
            6                                                                                                                                                                                                                                  -                                                                                                                                                                                                                          %         ,                                                                                                                                                                                                                               ,                                                                                                  	                                                                                                                         )          	    ,                   "                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                 -                  	                                                                                                                                                                                                         ,                                                                                                 

                                                                                                                     
         ,                                                                                                	                                                                                                                                           ,                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                 ,                                                                                                                                              
                                                         #                                ,                         	                                                                                                                 	                                                                                                  ,                                    
                                                                                                                                                           
                                       ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                           .               
                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                           ,          2                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                	        -                                                                                                                                                                                                                                         .                                                                                                                                                                                                                         ,                                                                                                                                    	                                                                                                  ,                                                                                                                                                                                                                                         -                                 #                                                                                                                                                                                                   /                          
                                                                                                                                                           	                                      ,                                                                                                                                     	                                                                                         -                                                                                                                                                                                                                  .                                                                                                                                                                                                                               ,                                  	                                                                                                                                                                         		                -                                                                                                                                                                                                                               .                                                                                                                                                                                                                         -                                                                                                                                                                                                                              -                                                                                                                                                                                                                 
       ,        
                                                                                                                                                                                                                   -                                                                                                                                                                                                                             .         
                                                                                                                                                                                                                1                                                                                                                                                                                                      ,                                                                                                                                                                                                                                 .                                                                                                                                                                                                                        .                                                                                                                                                                                                                     .                                                                                                                                                                                                                   -                                	                                                       
 	                                                                                                                                        .                                                                                                                                                                                                                     0                                                                                                                                                                                                                    .                                                                                                                                                                                                                                	     .                                                                                     	 	                                                                                                                        .                                                                                                                                                                                                                       .    
                
                                                                                                                                                                                                        ,                                                                                                                                                                                                                                          1                                                                                                                                                                                                  .                                                                                     	
                                                                                                                                  -                                                                                                                                                                                                                      /                                     	                                                                                                                                                                                         -                                                                                    
                                                                                                                      .                                                                                                                                                                                                            /                                                                                                                                                                                                                        0                                                                                                                                                                                                         2                                                                                                                                                                                                
/                                                                                                                          	                                                                       	.                                                                                                                                                                                                                  -                                                                                                                                     	                                                                                                 1                                                                                                                                                                                                         /                                                                                                                                                                                 
                         	        /                	                                                                                                                	                                                                                    .                                                                                                                                                                                                                              3                                                                                                                                                                                                       
.                                                                                                                                                                                                                $              -                                                                                                                                                                                                                       .                                                                                                                                                                                                                               .                                                                                                                                                                                                                         	-                                                                                                                                                                                                                     -                                                                                                                                                                                                                                          1                                                                                                                                                                                                   
    0               	                                                                                                                                                                                                      0                                                                                                                                                                                                       -                                                                                                                                  
                                                                                             -                                  
                                                                                                                                                                                          -       
                                                                                                                                                                                                                        .                                                                                                                                                                                                         
-                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                 .                                                                                                                                                                                                           	            0                                                                                                                                                                                                           0                                                                                                                                                                                                                      
    0                                                                                                                                                                                                  -    	                                                                                                                                                                                                                 -                                                                                                                                                                                           
/                                                                                                                                                                                                           	                 ,                                   	                                                                                                                                                                                  ,                                    
                                                       	                                                                                                                                   0                                                                                                                                                                                                      ,              	                                                                                                                                                                                                       .                                                                                                                                                                                                                                      .                                                                                                                                                                                                                   
,                                                                                                                                                                                                                   .                	     	                                                                                                                                                                                                        ,                                                                                                                                                                                                                                         1                                                                                                                                                                                                     -                                                                                      	                                                                                                                                  .                                                                                                                                                                                                                   0                                                                                                                                                                                                                        2                                                                                                                                                                                                   1                                                                                                                                                                                                          1                                                                                                                                                                                         
                         /                                                                                                                                                                                                             3                                                                                                                                                                                                /                                                                                                                                                                                                             .                                                                                           
                                                                                                                           ,                     
                                                                                                                                                                                                               3                                                                                                                                                                                                          0                                                                                                                                                                                                                    -                                                                                                                                                                                                           .                                                                                                                                                                                                                     /                                                                                                                                                                                                 .                                                                                                                                                                                                              #                ,      	                                                                                                                                                                                                                    .                                                                                                                                                                                                	                         
     .              	                                                                                                                                                                                                  /                                                                                                                                                                                                                          -     	                	              	                                                                                                                                                                                                     /                                                                                                                                                                                                            .                                                                                                                                                                                                                 .                                                                                                                                                                                                                               (      .                                                                                                                                                                                                                      -                                                                                                                                                                                                      	                   ,                                                                                          	                                                                                                                                .                     	                                                                                                                                                                                      
              /           
                                                                                                                                                                                                                      /                                                                                                                                                                                                                 
   .                                                                                                                                                                                                                0                                                                                                                                                                                                      
              -                                                                                                                                                                                                                            
      /                                                                                                                                                                                                            0                                                                                                                                                                                                      
/          	                                                                                                                                                                                                      "              -                                                                                                                                                                                                                           -                                                                                                                                                                                                                    .                                                                                                                                                                                                                                   .                                                                                                                                                                                                          	        /   	   	                                                                                                                                                                                                               -                                                                                                                                                                                                                                -                                                                                                                                                                                                           0                                                                                                                                                                                                             .  
                                                                                                                                                                                                                      0                                                                                                                                                                                                   /                                                                                                                           

                                                                                          .                                                                                              
                                                                                                                          .    
                    
   
                                                                                                                                                                                          0                                                                                                                                                                                                           2                                                                                                                                                                                                              1                                                                                                                                                                                                                      0                                                                                                                                                                                                                         1                                                                                                                                                                                                             	0                                                                                                                                                                                                  	.                                                                                                                                                                               
                               /                                                                                                                                                                                                           	/                                                                                                                                                                                                              1                                                                                                                                                                                                       .                                                                                                                                                                                                                           -                                                                                                                                                                                                                               .                                                                                                                                                                                                       
                  
     .                                                                                                                                                                                                         	3                                                                                                                                                                                                             /     	                                                                                                                                                                                                                     0                                                                                                                                                                                                   
            .                                                                                                                                                                                                                  ,                                                                                                                                                                                                                     .                                                                                                                                                                                                      /                                                                                                                                                                                                         	           .                                                                                                                                                                                                            	     -                
                                                                                                                                                                                                    !          .                  	                                                                                                                                                                                                            .                                                                                                                                                                                                                        -                                                                                                                                                                                                                      .                                                                                                                                                                                                               	    
-                    
                                                                                                                                                                                                               .                                                                                                                                                                                                             
         -                                                                                                                                                                                                                     2                                                                                                                                                                                                              -                                                                                                                                                                                                                             /                                                                                                                                                                                                               0                                                                                                                                                                                                       /                                                                                                                                                                                                                    -    	                                                                                                                                                                                                                           ,                                                                                                                                                                                                                        -                                                                                        
                                                                                                                                     -                                 	                                                                                                                                                                                           /                                                                                                                                                                                                             .                                                                                                                                                                                                                   
          .                                                                                                                                                                                                                     -                                                                                                                                                                                                           	         -                                                                                                                                                                                                                          /                                                                                                                                                                                                            .            	                                                                                                                                                                                                    -                                                                                            
                                                                                                                            /                                                                                                                                                                                                               .                                                                                                                                                                                                                1                                                                                                                                                                                                             0                                                                                                                                                                                                          -                                                                                                	                                                                                                                                  .                                                                                                                                                                                 	                                0                                                                                                                                                                                                         .                                                                                                                                	       
                                                                                     0                                                                                                                                                                                                         	       0                                                                                                                                                                                                          3                                                                                                                                                                                                  /                                                                                                                                                                                           
                         	    .             
                                                                                                                                                                                                                 .       	        	                                                                                                                                                                                                          1                                                                                                                                                                                                                   1                                                                                                                                                                                                     
         0                                                                                                                                                                                                                        -                                                                                                                                                                                                   	             /                                                                                                                                                                                                                     .                                                                                
                                                                                                                             /       
                                                                                                                                                                                                   .                                                                                                                                                                                                             	       -                                                                                                                                                                                                                  	.                 	                                                                                                                                                                                                 
          	      .                                                                                                                                                                                                                         .                              	                                                                                                                                                                                                .                                                                                                                                                                                                                       -                                                                                                                                                                                                                            -                 	                                                                                                                                                                                                                  /                                                                                                                                                                                                                  -                                                                                                                                                                                                                /                                                                                                                                                                                                                     0                   
                                                                                                                                                                                                   	      	    /                                                                                                                                                                                                         0                                                                                                                                                                                                        .                                                                                                                                                                                                                               -                                                                                                                                                                                                                             .                                                                                                                                                                                                           	         -                                                                                                                                                                                                                              /                                                                                                                                                                                                              .                                                                                                                                                                                                                   /                                                                                                                                                                                                               	               1                                                                                     
 
                                                                                                                           /                                                                                                                                                                                                  
             .         
         	           	                                                                                                                                                                                            /                                                                                                                                                                                                        ,                                                                                                                                                                                                                          .                                                                                         

                                                                                                                          -                           	                                                                                                                                                                                        .                                                                                                                                                                                                          .                                                                                                                                                                                                             
0                                                                                                                                                                                                              /                                      	                                                                                                                                                                                           2                                                                                                                                                                                                                 	0                                                                                                                                                                                                -                                                                                                                              
                                                                                       /                                                                                                                                                                                                        	          0                                                                                                                                                                                                        /                                                                                                                                                                                                       	.                                                                                                                                                                                        
                              .                                                                                                                                                                                                                               1                      	                                                                                                                                                                                                            0                                                                                                                                                                                                          0                                                                                 	                                                                                                                           -      	                                                                                                                                                                                                                            0                                                                                                                                                                                                                /                                                                                                                                                                                                                   -                                                                                                                                                                                                                /       
                                                                                                                                                                                                          0                                                                                                                                                                                                                   1                                                                                                                                                                                                                    /                                                                                                                                                                                                                          .                                                                                                                                                                                                              .                                                                                                                                                                                                                                 -                                                                                                                                                                                                                           .                                                                                                                                                                                                                         -                                                                                                                                                                                                                           .                                                                                                                                                                                                                                         -                                                                                                                                                                                                                
       /                                                                                                                                                                                                                     	-                                                                                                                                                                                                                      
        /            	                                                                                                                                                                                                      .                                                                                                                                                                                                                         .                                                                                                	                                                                                                                      '             .                                                                                                                                                                                                                    ,                                      6   	                                                                                                                                                                                              /                                 	                                                                                                                                                                                           ,                                                                                                                                                                                                 	                              -                                                                                                                                                                                                                   0                                                                                                                                                                                                                     -                                                                                                                                                                                                             0          	                                                                                                                                                                                              
         .                                                                                                                                                                                                              -                                                                                                                                                                                                                               3                                                                                                                                                                                                        1                                                                                                                                                                                                  
                .                                                                                                                                                                                                                   /                                                                                                                                                                                                         /                                                                                                                                                                                                                  /                                                                                                                                                                                                                 /                                                                                                                                                                                         	                                 /                                                                                                                                                                                                       0                                                                                                                                                                                                    
.                                                                                                                                                                                                                  .                                                                                                                                                                                                                       -                                                                                                                                                                                                                          2                                                                                                                                                                                                      	/                                                                                                                                                                                                                         .            	                                                                                                                                                                                                    /                                                                                                                                                                                                              	                           1                                                                                                                                                                                                              
0                
                                                                                                                                                                                                       .                                                                                                                                                                                                                         -                                                                                                                                                                                                                         0                 
                                                                                                                                                                                               /                                                                                                                                                                                                                        /                	                                                                                                                                                                                                  0                                                                                                                                                                                                                 
      -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                    9   
       .              	                                                                                                                   
	                                                                                     -                                                                                                                                                                                                                                   -                                                                                                                                                                                                                                   .                                                                                                                                                                                                                  
        -        	                                                                                                                                                                                                  	        	     .                                                                                                                                                                                                                           /                                                                                                                                                                                                       
           /                                                                                                                                                                                                          	              
   /                                                                                                                                                                                                                    0                                                                                                                                  	
                                                                                       .                                                                                                                                                                                                                -                                                                                                                                                                                                                              ;              .                                                                                                                                                                                                                    .                                                                                                                                                                                                  .                                                                                                                                                                                                              ,                                                                                                                                                                                   	                                .                                                                                    
                                                                                                                                    .                                                                                                                                                                                                                                   -                                                                                                                                                                                                          	              /                          	                                                                                                                                                                                     -                     
                                                                                                                                                                                                              /                                                                                                                                                                                                               '                ,     
                                                                                                                                                                                                        	
                1                           
                                                                                                                                                                              -                                                                                                                                                                                                                  .                                                                                                                                                                                                      	            /                                                                                      
                                                                                                                                 .                                                                                                                                                                                                                               .                                                                                                                                                                                                             2                                                                                                                                                                                                           	0                                                                                                                                  
                                                                            /                                                                                                                                                                                                             2                                                                                                                                                                            	                              /         	                                                                                                                                                                                                              "       ,                 	                                                                                                                                                                                                         1                                                                                                                              
                                                                                         -          
                                                                                                                                                                                                          -                                                                                                                                                                                                               
                  
     /                                                                                                                                                                                                                              	 .                                                                                                                                                                                                               ,      
            
                                                                                                                                                                                                             0                                                                                                                                                                                                              -                                                                                                                                                                                                                   ,                                                                                                                                                                                                                         .                                                                                                                                                                                                             .                                                                                                                                                                                                           
     .                                                                                                                                                                                                                            .                                                                                                                                                                                                                          +          -                                                                                                                                                                                                                 .                                                                                                                                                                                                                                 .                                                                                                                                                                                                                
     
          /                                                                                                                                                                                                                        1                                                                                                                                                                                                                             ,                                                                                                                                                                                                                         ,                                                                                                                                                                                                                      
  0                                                                                                                                                                                                               
    
       /                                                                                                                                                                                                                  .                                                                                                                                                                                                                       /                                                                                                                                                                                                            -                                                                                                                                                                                                                           ,           
     .                             
                                                                                                                                                                                       /                                                                                                                                                                                                     -                         	                                                                                                                                                                                   /                                                                                                                                                                                                                   .                                                                                                                                                                                                      /                  	                                                                                                                                                                                           	                        /                                                                                                                                                                                                                          
 .                              
                                                                                                                                                                               .                                                                                                                                                                                                                                      .                                                                                                                                                                                                             "               -                                                                                        	                                                                                                                               2                                                                                                                                                                                                         .      	             	                                                                                                                                                                                                      /                                                                                      
                                                                                                                              0                                                                                                                                                                                                                  .                                                                                                                                                                                                                                   0                              	                                                                                                                                                                                     0                                                                                                                                                                                                         0                                                                                                                            	                                                                        .                                                                                                                                                                                                          /                                                                                                                                                                                                    0                                                                                                                                                                                                                          -                                                                                                                                                                                                           -                                                                                                                                                                                                                            ,          	     	       	                                                                                                             	                                                                                                -                                                                                                                                                                                                                     	          
     .                                                                                                                                                                                                                  	       	        /                                                                                                                                                                                                      -  	      	                                                                                                                                                                                                                     /                                                                                                                                                                                                              -                                                                                                                                                                                                                   -                               
   
                                                                                                                                                                                                  2                                                                                                                                                                                                                /                                                                                                                                                                                                                          -                                                                                                                                                                                                                         -                                                                                                                                                                                                      	                         .  
     /                  
                                                                                                                                                                                                     -                                                                                                                                                                                                                               -                                                                                                                                                                                                                                    .                                                                                                                                                                                                                          .           
                                                                                                                                                                                                           ,                                                                                                                                                                                                                         ,                                                                                                                                                                                                                      /                                                                                                                                                                                                               
          /             	                                                                                                                                                                                                     /                                                                                                                                                                                                 	              .                                                                                                                                                                                                           ,                                                                                                                                                                                                                        	       @                   .                                                                                                                                                                                                                   .                                                                                                                                                                                                           -                                                                                                                                                                                                                -                                                                                                                                                                                                                 ,                                                                                                                                                                                                               /                                                                                                                                                                                                                     	           .                                                                                                                                                                                                                    .                                                                                                                                                                                                              ,   
                                                                                                                                                                                                                                   .                                                                                                                                                                                                                              -   	             
                                                                                                                                                                                              	                 2                                                                                                                                                                                                                -                                                                                                                                                                                                                 -                                                                                                                                                                                                              -                               	                                                                                                                                                                                             -                                                                                                                                                                                                                              .                                                                                   
 
                                                                                                                                    -                                                                                                                                                                              	                                /                                                                                                                                                                                     
                             	.                                                                                                                                                                              
                               
/                                                                                                                                                                                                          1                                                                                                                                                                                                                          -                                                                                                                                                                                	   
                         0                                                                                                                                    	                                                                                     ,                     
                                                                                                                                                                                                            /                                                                                                                                                                                                               
          	     /                                                                                                                                                                                                         
                1                                                                                                                         
                                                                                        ,        
                                                                                                                                                                                                                       /                                                                                                                                                                                                        .                                                                                                                                                                                                                   -                                                                                                                                                                                                                           -                                                                                                                                                                                                            	/                                                                                                                                                                                                                          ,                                      
                                                                                                   
                                                                                                 -                                                                                                                                                                                                    	            	            
    ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                   1     
     ,                                                                                                                                                                                               
                                 -                                                                                                                                                                                                                       $        ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                             "         
   -                     
                                                                                                                                                                                                     -                                                                                                                                                                                                                                       ,                          
                                                                                                                                                                                                         -                                                                                               	                                                                                                                           -                  
                                                                                                                                                                                                                 .                                                                                                                                                                                                               ,                                                                                                                                                                                                                           ,                                      	                                                                                                                                                                                            ,                                                                                                                                                                                                                                .                                                                                                                                                                                                                           ,                                                                                                                                                                                                                        -                                                                                                                                                                                                                   	               ,                   .                                                                                                                                                                                                                               /                                                                                                                                                                                                                                   
   -                                                                                                                                                                                                           ,                                                                                                                                                                                                                            -         
       ,                                                                                          	                                                                                                                                        	/                                                                                                                                                                                                                      0                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                       ,                                    
                                                                                                                                                                                              /                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                    /                                                                                                                                                                                                               
        1                                                                                                                                                                                                                       .                                                                                                                                                                                                                                	      -                                                                                                                                                                                                                                             -                                                                                                                                                                                                                                 0             
                                                                                                                                                                                                 ,                                                                                             
                                                                                                                                       -                                                                                                                                                                                                                                      -                                                                                                                                                                                                                                 /                                                                                                                                                                                                               /                                                                                                                                                                                                                            ,                                                                                                                                       .                                                                                                  1                                                                                                                                                                                                                             -                                                                                                                                                                                                                          -                                     	                                                                                                                                                                                    %   
     ,                                    
                                                                                                                                                                                            -                                                                                                                                                                                                                                -                                                                                                                                                                                                                 
           -                                                                                                                                                                                                                             /          -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                        -                                                                                                                                                                                                           	   
          ,                                                                                                       	                                                                                                                   	       !                  .                       
                                                                                                                                                                                                         ,                                                                                                                                                                                                                                                 .                                                                                                                                                                                                                       	        ,                                                                                                                                                                                                                          ,                                
                                                          	                                                                                                                                    .                                                                                                                                                                                                                           -                      	                                                                                                                                                                                                        ,                                                                                                                                                                                                                          	         ,                                                                                                                                 	                                                    	                                -                                                                                                                                                                                                                            -                                                                                                                                                                                                                    -           	                                                                                                                                                                                                                   -                                                                                                                                                                                                                                     ,                                                                                                                                                                                                  	                               /                                                                                                                                                                                                      	        ,                                                                                                                                                                                                                         #           	    -                                                                                                                                  	                                                                                          ,                                                                                                                                                                                                                                   
      ,                             
                                                                                                                                                                                              -                                                                                                    	                                                                                                                        
             ,                                                                                                      
                                                                                                                                             ,                                                                                         
                                                                                                                                              ,                                                                                                                                                                                                               
                ,                                                                                                                                                                                                           
                             
       ,                                                                                                                                                                                                                                          "        -                 
                                                                                                                       #                                                                                                     ,                                                                                                   	                                         	                                                      	                                     ,                                                                                                                                                                                                                              &             ,                                                                                                                                                                                                                                    
,                                                                                                     	                                                                                                                                        -                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                        -                                                                                                                                                                                                                                            .                                                                                           	                                                                                                                                    .                                                                                                                                                                                                                            0                                                                                                                                                                                                                        -                                                                                                                                 $                                                                                       -                                                                                                                                                                                                                         ,                                                                                                                                                                                                                              -                                                                                                                                                                                                                           /                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                  8          -                                                                                                                                  	                                                                                           .                                                                                                                                                                                                                                   $         ,                   #       	                                                                                                                                                                                                       	           -                                                                                                                                                                                                                                   -                                                                                                                                                                                                                 	                 ,                                                                                                                                                                                                                                            ,           %              	                                                                                                                                                                                                       	           -          
                                                                                                                                                                                                                         -           	            	                                                                                                                                                                                                             ,                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                 -                                                                                                     	                                                                                                                   )
                ,                                                                                                                                                                                                                             ,                                       C                                                                                                                                                                                                 -         	                                                                                                                                                                                                                     .                                                                                                                                                                                  	                                -                                                                                                                                                                                        	                                    -                                                                                                                                                                                                          	                             4   	        -        
  '                                                                                                                                                                                                                             ,            	                                                                                                                                                                                                                     -                                                                                                                                                                                                                          -                                                                                              	                                                                                                                             $                   ,                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                              -                 	                                                                                                                                                                                                        ,                                                                                                      
                                                                                                                           $                  ,                                                                                                   '                                                                                                                                       ,                                                                                                                                                                                                                               0                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                    
            	     ,                                                                                                                                                                                                                 %                                /                   	                                                                                                                                                                                                             ,                                                                                                                                        %                                                            	                                        ,                                                                                                                                                                                                          	                            #          .                                                                                                                                                                                                                             ,                                                                                                                                                                                                     
                             -                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                        /                  )                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                    4           -                       	                                                                                                                                                                                                         	     ,                                                                                                                                                                                                                                        .                                                                                                                                                                                                                          /                                                                                                                                                                                                                -                                	                                                                                                                                                                                           ,                                                                                                                                                                                                                                    ,          
                                                                                                                                                                                                                     -                                                                                                                                                                                                                            	              -                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                              /             ,                 ,                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                  -                #                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                 
      .         ,            "                                                                                                                                                                                                                                      -                                                                                                                                                                                                                                      ,                     "                                                                                                                                                                                                                               -                                                                                                                                                                                                                             ,       
                                                                                                                                                                                                                         ,                                                                                                                                                                                                                           6              ,                                                                                                                                                                                                                                   .                                                                                                                                                                                                                             ,                                 
                                                                                                                                                          
                                  
,         	                           >                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                         -         @                                                                                                                                                                                                                                      .                                                                                                                                                                                                                           ,                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                                   0                                                                                                                                                                                                                        -       	                                                                                                                                                                                                              ,                                    	                                                                                                                                                                                                      ,                                                                                                                                                                                                                                         -                                                                                                                                          
                                                                                              ,                              !                                                                                                                                                                                                  ,                                                                                                                                                 )                                                                                                     ,                                                                                                                                                   	                                                            5                                      ,                                                                                                                                           	                                                           %                                        ,                                                                                                                                          5                                                            	                                         -                                                                                                                                                                                                                               ,                                                                                                                                                                                                                                                  -                                                                                                                                                                                                                             .           	
                                                                                                                     	                                                                                ,                                                                                                                                                                                                                              -                                                                                                                                                                                                                               /                 	                                                                                                              
                                                                                        -            	                                                                                                                                                                                                            -                                                                                                                                                                                                                             -                                                                                                                                                                                                               ,      
   	                                                                                                                                                                                                                                    ,       	                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                            	    ,                    
                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                       -                                                                                                                                                                                                                                      -                                                                                                                                                                                                                              .                    ,           $                                                                                                                                                                                                                              -                                                                                                                                                                                                                                     ,          
                                                                                                                                                                                                              	                 ,                                                                                                                                                                                                                                               ,                                       	                                                                                                                                                                                                -                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                        ,                                                                                                   	                                                                                                                           -                                                                                                                                                                                                                                    ,                	                                                                                                                                                                                                          7             -                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                  ,                                       $                                                                                                                                                                                                         ,                                         
                                                          	                                                                                                                                      ,                 	                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                              ,             '                                                                                                                                                                                                                                            -                                                                                                                                                                                                                                
    ,                  
                                                                                                                                                                                                        ,                   
       
                                                                                                                                                                                                                     ,                  
                                                                                                                      	                                                                                                -                                                                                                                                                                                                                         
     ,      	                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                     -                                     &   
                                                                                                                                                                                                   ,           	                           	                                                                                                                                                                                                            ,                                                                                                                                                                                                                                  ,                        
                                                                                                                                                                                                                -                                                                                                                                                                                                                                  ,                                                                                                                                    
                                                                                                      ,                  	                                                                                                                                                                                                                           -                                                                                                                                                                                                                        	           -                   
                                                                                                                                                                                                              ,                                                                                                                                                                                                                                   ,             <                                                                                                                                                                                                                                           -                                                                                                                                                                                                                               ,       	                                                                                                                                                                                                                       ,                                                                                             	                                                                                                                                       ,                     .                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                	              ,                      	             	                                                                                                                                                                                                   -                                                                                                                                                                                            	                               ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                            "        -                                                                                                                                                                                                                           -                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                      	              &              ,                                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                             &       ,                                                                                                                                                                                                                                              -                                                                                                                                                                                                                                     '              ,                                                                                                                                                                                                                                       -                                                                                             	                                                                                                                                      ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                               G               ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                             -                                                                                                                                                                                                                        	            .                                                                                                                                                                                                                      /             -                 )                                                                                                                                                                                                                      -               	                                                                                                                                                                                                                  .                  ,      	                                                                                                                                                                                                                       .                                                                                                                                                                                                            
           ,                	                                                                                                                                                                                                                             ,                                                                                                                                                                                                                           +                 .                                                                                                                                                                                                                                 -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                    9            
,                                                                                                                                                                                                                                               .                                  	                                                                                                                                                                                           0                                       .                                                           
                                                                                                                                              ,                                                                                                                                                                                                                             	               ,                                                                                                                                                                                                                               	        -                                                                                                                                                                                                                          -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                             -              /                                                                                                                                                                                                                           ,              	                                                                                                                       	                                                                                           -                                                                                                                                  	
                                                                                              .                                                                                                                                                                                                                                        -                                                                                                                                                                                                                                       	     	.                                                                                                                                                                                                                            ,               &                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                            
    	   .                 	                                                                                                                                                                                           
                  ,          2                                                                                                                                                                                                                                   -                                                                                                                                                                                                                   ,                                                                                                                                                                                                                         ,                                                                                                                                                                                                	                                    .                 	#                                                                                                                                                                                                                   ,                                                                                                                                                                                                                               &        /                                                                                                                                                                                          	                                  -                                                                                                                                                                                                                      	               	   .                                                                                                                                                                                                                        ,                                                                                                                                                                                                                             	    ,                                                                                                                                                                                                                            .                                                                                                                                                                                                                          
   /                                                                                                                                                                                                                          ,                  	                                                                                                                    	                                                                                        ,                                                                                                                                                                                                                     ,                                                                                                                                                                                                                     +               /                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                 -                                                                                                                                                                                                                      -                                                                                                                                                                                                                       /                                                                                                                              	                                                                                             /                                                                                                                                                                                                                     .   
                                                                                                                                                                                                                             -                                                                                                                                                                                             	                               .                                                                                                                                                                                                                    ,                                                                                                                                                                                                               
              .                                                                                                                                                                                                                -                                                                                                                                                                                                                      .                                                                                                                                                                                                           ,        
                                                                                                                             
                                                                                                  ,                                    	                                                       	                                                                                                                    	              /                                                                                                                               	                                                                                      /                                                                                                                                                                                                                                 -          	                                                                                                                                                                                                             -                                                                                                                                                                                                                             /                                                                                                                                                                                                                          -                                                                                                                                                                                     	                                     -                                                                                                                                                                                                                               0            "             
                                                                                                                                                                                                              2                                                                                                                                                                                               	                       	   .                 

                                                                                                              
                                                                                         -                                                                                                                                 
                                                                                       .                                                                                                                                                                                                                               1                                                                                          	                                                                                                                           	-                                                                                                                                                                                                                         .                                                                                                                                                                                                                       -                                                                                                                                                                                                                      /                 	                                                                                                            	                                                                                    /                                      
                                                                                                                                                                                 ,                                                                                                                                                                                                                     
    -                  
	                                                                                                                     	                                                                                  .                                                                                                                                                                                                                           #        ,                                                                                                                                                                                                                                           
,                                                                                                                                                                                                                              $	                0                                                                                                                                                                                                                      ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                               -                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                ,                                                                                                                                                                                                                     -                                                                                                                                                                                                                             #              ,                                                                                                                                                                                                                                    .                                                                                                                                                                                                                                   .                                                                                                                                                                                                                     -                                                                                                                                                                                                                             ,            	                                                                                                                                                                                                                       ,                                                                                                                                                                                                                             	       +                     ,                 $                                                                                                                                                                                                                         /                                                                                                                                                                                                                      -                                                                                                                                                                                                                                          -                                                                                                   	                                                                                                                             ?                    -                                                                                                                                                                                                                                      .                                                                                                                                                                                                                     -                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                           
      -                                                                                           #                                                                                                                                         ,                                                                                                                                                                                                                               /                                                                                         
                                                                                                                                         ,                                                                                                                                                                                                                                        
   
   .                                                                                                                                                                                                                                 .                                                                                                                                                                                      
                             -                                                                                               
                                         -                                                                                               ,                                                                                                                                                                                                                                      -           .                 
                                                                                                                                                                                                               -                                                                                                                                                                                                                           ,                                                                                                                                                                                                                        ,                                                                                                                                                                                                                           
             ,            -                      
                                                                                                                                                                                                        /                                                                                                                                                                                                                 ,          %                                                                                                                                                                                                                                ,                                                                                            
                                                                                                                                  -                                                                                                                                                                                                                          ,                                                                                            
                                                                                                                                ,                                                                                                                                                                                                                   
              ,                            
         
                                                       	                                                                                                                                        ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                     
        ,                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                               .                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                       	             ,                  (                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                          #             -            
                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                        	      -                                                                                        	                                                                                                                                -                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                              ,                          
                                                                                                                                                                                                            ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                               .                                                                                                                                                                                                                    	      ,                                                                                                                                                                                                                                    .                                                                                                                                                                                                                           #     
   ,                                                                                                                                                                                                                                           0                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                       -                                   	                                                                                                                                                                                                       ,                                                                                                                                                                                                                                     .                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                	             ,                                                                                                                                                                                                                                    
   ,                                      %                                                                                                                                                                                                               .                                                                                                                                                                                                               ,                                                                                                                                                                                                                               !        ,                                                                                                                                                                                                                %                          
             ,                                                                                                                                             ,                                                                                                .                                                                                                                                     	                                                                                             ,                                                                                                                                                                                                                                          +             ,                                                                                                                                                                                                                                       -                                
                                                                                                                                                         
                                     -                                                                                                                                                                                                                 .                                                                                                                                                                                                                               +            ,      	                                 	                                                                                                                                                                                                      .                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                      	              ,                                                                                                                                                                                                   
                         .                                                                                                                                                                                                                                ,                
                                                                                                                                                                                                                      ,                                                                                                                                                                                            
                               /              
                                                                                                                                                                                                -                                                                                                                                                                                                                      
                 -                                                                                                                                                                                                                          /                                                                                                                                                                                                                              /                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                   	   /                                                                                                                                                                                                                     .                                                                                                                                                                                        	                           /     
               	                                                                                                                                                                                                          ,                                                                                                                                                                                                                                        0     	                                                                                                                                                                                                                -                                                                                                                                                                                                                                  /                                                                                                                                                                                                                ,                                                                                                                                                                                                                   	                 .                                                                                                                                                                                                                -                                                                                                                                                                                                               -                                                                                                                                                                                                                     0                                                                                                                                                                                                               -               	                                                                                                                                                                                                               -                                                                                                                                                                                                                       
            .                                                                                                                                                                                                               	0                                                                                                                                                                                                                ,  	               
                                                                                                                                                                                                               .                                                                                               	                                                                                                               #                -              !                                                                                                                                                                                                                   -                                                                                                                                                                                                                        /                                                                                                                                                                                                                     .                                                                                      
                                                                                                                         .                                                                                                                                                                                                                       .                                                                                                                                                                                                                   2                                                                                                                                                                                                                     0                                                                                                                                                                                                   1                                                                                                                                                                                                                0                                                                                                                                                                                                                  0                                                                                                                                                                                                                   .                                                                                                                                                                                               
                               	    ,                                                                                                                                                                                                                             /                                  	                                                                                                                                                                             
      /                                                                                                                                                                                                                 .                                                                                                                                                                                                                                    .                                                                                                                                                                                                   
          -                                                                                                                                                                                                        .                                                                                                                                                                                                                      0                                                                                                                                   	                                                                                  .                                                                                                                                                                                                                
.                                 
                                                        	                                                                                                                   
                ,
  
                                                                                                                                                                                                                                 /                                                                                                                                                                                                      0                                                                                                                                                                                                                  ,                                                                                                                                                                                                                           2       -                
                                                                                                                                                                           	                             .                                                                                                                                                                                                                            ,                                                                                                                                                                                                                          /                                                                                                                                                                                                                         -      	                                                                                                                                                                                                                               ,                                                                                                                                                                                                                   
             .                                                                                                                                                                                                                        -                                                                                                                                                                                                                 	           ,                    
                                                                                                                                                                                                             -                                                                                    
                                                                                                                               .                                                                                                                                                                                                            .                                                                                                                                                                                                                 
       -                .                             	                                                                                                                                                                                         0                                                                                     
                                                                                                                                ,                                                                                      
                                                                                                                                     ,                                                                                                                                 	                                                                                          0                                                                                                                                                                                                                /                      
                                                                                                                                                                                                               ,                                                                                                                                                                                                                        	  -                                   	                                                                                                                                                                                -           
                                                                                                                                                                                                               .                   	                                                                                                                                                                                                          ,                                                                                          	                                                                                                                   
           0                                 
                                                                                                                                                                                      .                                                                                                                                                                                                                              /                                                                                                                                                                                                                   
0                                                                                                                                                                                                             .                                                                                              
                                                                                                              
             0                                                                                                                                                                                                             
         0                                                                                                                                                                                                      
1                                                                                                                                                                                                              ,                                                                                                                                                                                                           .                                                                                                                                                                                                             .                                                                                                                                                                                                                            -                                                                                                                                                                                     	                             /                                                                                                                                                                                                                            -                                                                                                                                                                                                                        .         	     
     	                                                                                                                                                                                                               -                                                                                                                                                                                                                   0                                                                                                                                                                                                     .                                                                                                                                                                                                                            /                                                                                                                                                                                                                      -                   
                                                                                                                     
                                                                                 -                                                                                                                                                                                                                        /        	                                                                                                                                                                                                              0                                                                                                                                                                                                            /                                                                                                                                                                                                              ,                                                                                                                                                                                                                         )    
  .                                                                                                                                      	                                                                                  -                                                                                                                                                                                                                                .                                                                                                                                                                                                                     -                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                               .                                                                                                                                                                                                                    
    0                                                                                                                                                                                                                 ,                                                                                                                                                                                                                            -                                                                                                                                                                                                                               .                                                                                                                                                                                                                  .                                                                                                                                                                                                            -                                                                                                                                                                                                                         *               .                                                                                                                                                                                                                           /                                                                                                                                                                                                                   /                                                                                                                                                                                                                  .                                                                                                                                                                                                                 -                                                                                                                                                                                                -                                                                                                                                                                                                                                -                                                                                                                                                                                                                -          
                                                                                                                                                                                                     .   	           
                                                                                                                                                                                                        /                                                                                                                                                                                                                              /                                                                                                                                                                                                           0                                                                                                                                                                                                                  /   	  	                                                                                                                                                                                                            1                                                                                       
                                                                                                                          0                                                                                                                                                                                                           /                                                                                                                                                                                                    1                                                                                                                                                                                                                     1                                                                                                                                                                                                      .                                                                                                                                                                                              
0                                                                                                                                                                                                    
.                                                                                                                                                                                                                  .    	       	        	                                                                                                                                                                                                     -                                                                                                                                                                                                          /                                                                                                                                                                                                                      .        	                                                                                                                                                                                                              -                                                                                                                                                                                                                                 3                                                                                                                                                                                                                    	0                                                                                                                                                                                                              /                    	                                                                                                                                                                                                -                                                                                                                                                                                                                       -                                                                                                                                     	                                                                                 .    
                                                                                                                                                                                            
             .                                                                                                                                                                                                             /                                  
                                                                                                                                                                             	       -                                                                                                                                                                                                                          	      ,                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                       	.                                                                                                                                                                                                                          -                                                                                                                                                                                                                              -                                                                                                                                                                                                                               .                                                                                                                                                                                                                     ,                                                                                                                                                                                                                         
                 -                                                                                                                                                                                                                   
         
,      	                                                                                                                                                                                                                          .                                                                                                                                                                                                                             -         
                          
                                                                                                                                                                                        -                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                               /                                                                                                                                                                                                                      -                                                                                                                                                                                                                                ,                                                                                                                                            	                                                         
                             -                         	                                                                                                        	                                                                                         -        	                                                                                                                                                                                                                      .                                                                                                                                                                                                                     
           .                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                   -                                                                                                                                                                                                                       !                   ,                  
                                                                                                                                                                                                             0                                                                                                                                                                                                                       ,               	                                                                                                                                                                                                          ,                                                                                                                                                                                                                                  
-                                                                                        
                                                                                                                                      	-                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                  -                                                                                                                                                                                                                             -                                                                                                                                                                                                                                
-                                                                                                                                            	                                                                                          -                                                                                                                                                                                                                .                 	                                                                                                                                                                                                       -                                                                                                                                	                                                                                               -                                                                                                                                                                                                                       -                    
                                                                                                                                                                                                                   -                                                                                                                                                                                                                           .          	      
                                                                                                                                                                                                            /                                                                                                                                                                                                                  -                                                                                           
                                                                                                                    	                ,                                                                                                                                                                                                                         ,                                                                                        
                                                                                                                                    -                               
                                                                                                                                                                                           ,                                                                                                                                                                                                                                      
-                                                                                                                                                                                                                           .                                                                                                                                                                                                                                     -                                                                                                                                                                                                                            $        ,                                                                                                                                                                                                                           -                                                                                                                                                                                                                   
           
    ,               	                                                                                                                                                                                                    ,                                                                                                                                                                                                                                     ,          	                                                                                                                                                                                                
                 ,                                                                                                                                                                                                                             "             -        	                                                                                                                                                                                                             -                                                                                                                                                                                                                       .            
                                                                                                                                                                                                                 
      .                                                                                                                                                                                                                              ,                                                                                                                                                                                                                               /                                                                                                                                                                                                               #                  -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                   /                                                                                                                                 	                                                                                     -                                                                                                                                                                                                                                ,                                                                                                                                             	                                                                                                     -                                                                                                                                                                                                                            
       .                                                                                                                                                                                                                     0                                                                                                                                                                                            
                  	         ,                                                                                                                                                                                                                        /                                                                                                                                                                                                               
                         ,                                                                                                                                 	                                                          
                           
.                                                                                                                                                                                                                         -       	                                                                                                                                                                                                                         -                                                                                                                                                                                                                        /                                                                                                                                                                                                                    
           -                                                                                                                                                                                                                                       ,                                  	                                                                                                                                                                                           -                                                                                                                                                                                           	                          ,                                                                                                                                                                                                        
                             ,                                                                                                                                                                                                                                              -                  	                                                                          
                                                                                                                                  .                                                                                                                                                                                                    
                           
      ,                                                                                                                                                                                                                              -                                                                                                                                                                                          	   	                    	        -                                                                                                                                                                                                                                -         	                                                                                                                                                                                                                      ,                                                                                                                                                                                                                            .                                                                                                                                                                                                               .                                                                                                                                                                                                                      ,                                                                                            
                                                                                                                         
       -                                                                                                                                                                                                                              -                                                                                              
	                                                                                                                                   	      ,     	                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                            -                
                                                                                                                                                                                                                     -              	                                                                                                              	                                                                                       -                                                                                                                                                                                                                                 -           	                                                                                                                                                                                                                  
     ,                                                                                                                                                                                                                                          .                                                                                                                                                                                                       
           .                                                                                                                                                                                                                   -                       	                                                                                                                                                                                                          -                                                                                                                                                                                                                                        .                                                                                                                                                                                                              	      ,                                                                                                 	                                                                                                                     	          .                                                                                                                                                                                                                                   -                                                                                                                                                                                                                          	          .                                                                                                                                                                                                              /                                                                                                                                                                                                                      	  ,                                                                                                                                     
                                                                                           ,                                                                                                                                            /                                                                                               /                                                                                                                                                                                                                 .                                                                                                                                                                                                             	       /                                                                                                                                                                                                                    .                                                                                                                                                                                                                   -               
                                                                                                                        	                                                                                              .                                                                                                                                                                                                                      
-                                                                                                                                                                                                                  -                                                                                                                                                                                                           -                                                                                                                                                                                                                                   ,                                                                                                $ 	                                                                                                                                           .                                                                                                                             
                                                                                     -                                                                                                                                                                                        
                                    ,                               '                                                                                                                                                                                                       ,                                                                                                                                                                                                       	   #                         	       .                                                                                                                                                                                                                   /                                                                                            
                                                                                                                              0                                                                                                                                                                                                                                /                                                                                                                                                                                                                                 /          
                                                                                                                                                                                                               /                                                                                                                                                                                                                 -                                                                                                                                                                                                                           -                                                                                                                                                                                                                              ,          	    
                                                                                                                                                                                                              1                                                                                        	                                                                                                                                /      	                                                                                                                                                                                                              -                                                                                                                                                                                                                                 .                                                                                                                                                                                                                           .                                                                                                                                                                                                                        -                                                                                                                                                                                                                                     -                                                                                                                                                                                                                            ,                                                                                                                                                                                                                   -                                                                                                                                                                                                              	           -          
                                                                                                                           	                                                                                             -             
                                                                                                                                                                                                            	   -         
                                                                                                                                                                                                        ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                       .                                                                                                                                                                                                                  	      -         	  	                                                                                                                                                                                                           ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                         -                                                                                                                                                                                                                            .                                                                                                                                                                                                               -                                                                                                                                                                                                                     
       ,                                                                                                                                                                                                                               -                                                                                                                                                                                               
                                	-               	                                                                                                                                                                                                                     -                                                                                                                                                                                                                            	      ,               	                                                                                                                                                                                                                     -                                                                                                                                                                                                                                                  -                                                                                                                                        	                                                                                          0                                                                                                                                                                                                                      -                                                                                                                                                                                                                          ,                                                                                                  	                                                                                                                             &                  ,                                                                                                                                                                                                                         .                                                                                                                                                                                                                          -                                                                                                                                                                                                                    -                                                                                                     
                                                                                                                      	           .                                                                                                                                                                                                                               
,                                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                           	                             	    ,                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                           -                                                                                                                                                                                                                 -                                                                                                                                                                                                                                     -           	                                                                                                                                                                                                                      .                                                                                                                                                                                                               	       ,                                                                                                                                                                                                                         ,                                                                                                                                                                                                                       3            ,            !                                                                                                                                                                                                                          /                                                                                                                                                                                                                      -                                                                                                                                                                                                                    -                                                                                                                                                                                                                     /                                                                                                                                                                                                                             /                                                                                                 

                                                                                                                   	          	   -                                                                                                                                                                                                                                .                                                                                                                                                                                                                             ,                                                                                                                                                                                                                            ,                                   	                                                                                                                                                                                           -                                                                                                                                                                                                                         ,                                                                                                                                                                                                                 	       -            	                                                                                                                                                                                                                        ,               	                                                                                                                                                                                                                 .           
                                                                                                                                                                                                                          	      -                                                                                              	                                                                                                                   ,                                                                                                                                                                                                                                         ,       	                                                                                                                                                                                                                  -                                                                                                                                                                                                                        
             	    ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                                   ,               	                                                                                                                	                                                                                  
     .                                                                                                                                                                                                                                   /                                                                                                                                                                                        
                            .                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                     ,                
                                                                                                                                                                                                                        	,                                                                                                                                                                                                                              &           	     ,                  -                                                                                                                                                                                                                            /                                                                                                                                                                                                                    -                                                                                                                                                                                                                             -                                                                                                                                                                                                             	                   ,                                                                                                                                                                                                                                     .                                                                                                                                                                                                                    -      	   	                                                                                                                                                                                                             ,                                                                                             
                                                                                                                     
              
,                                                                                                                                                                                                                       		           ,                                                                                                                                                                                                                                    -         
                                                                                                                                                                                                                               ,                                                                                                                                                                                                                          ,                                                                                                                                                                                                       
                          ,                                                                                                                                                                                                                                            .                                                                                                                                                                                             	                                     -                                                                                                                                                                                                	                                 .                                   	   	                                                                                                                                                                                          
-                                                                                                                                                                                        	                            ,                                                                                                                                                                                                                            -                                                                                                                                                                                                             	       
                  ,                                        
                                                                                                                                                                                                  -                                                                                                                                                                                               
               ,                                                                                                                                                                                                                  	               .                      	                                                                                                                                                                                                            ,             	                                                                                                                                                                                                            ,                                                                                                                                                                                                                                           /                                                                                                                                                                                                                              /                                                                                                                                                                                                             -                                                                                                                                                                                                                  /                                                                                                                                                                                                                   .                                                                                                                                                                                                                           -                                                                                                                                                                                                                                -                                                                                          	                                                                                                                               -            	                                                                                                                                                                                                       	                    /           
                                                                                                                                                                                                                 ,                  	                                                                                                                                                                                                           .          	       	                                                                                                                                                                                               /                                                                                                                                                                                                                                           .   
                                                                                                                                                                                                                           -                                                                                   	                                                                                                                       
              .                                                                                                                                                                                                                    /                                                                                                                                                                                                                   .          .                                                                                                                                                                                                                   -                                                                                                                                                                                                                /                                                                                                                                                                                                                     ,                                                                                                                                                                                    	                                     	-                                                                                          	                                                                                                                                 .                                                                                                                                                                                                                                  -                                      
                                                                                                                                                                                      /                                                                                                                                                                                                                   -    	         	                                                                                                                                                                                                                         ,                                                                                                                                                                                                                           /                                                                                                                                                                                                        
0                                                                                    	                                                                                                       	             -                           	                                                                                                                                                                                                  .                                                                                                                                                                                                                   	0                                                                                       
                                                                                                                            -                             
                                                                                                                                                                                    /                                                                                                                                                                                                                 1                                                                                                                                                                                                                    1                                                                                                                                                                                                      1                                                                                                                                                                              	                           	.                                                                                                                                                                                                                  -                                                                                                                                                                                                                          -                                                                                                                                                                                                    1                                                                                                                                                                                                                0            	                                                                                                                  
                                                                                          .                                                                                                                                                                                                       	                      .                                                                                                                                                                                                                     
/                                                                                                                                                                                          
               -                                                                                                                                                                                                                               .                                                                                                                                                                                                                            .                                                                                                                               	                                                                                     ,                                                                                        	                                                                                                                              ,                                                                                                                                                                                                                      .                                                                                                                                                                                                               
       .               
                                                                                                                                                                                                     .                                                                                                                                                                                          	                         	  ,                                                                                                                                      	 
                                                       	                            ,                                                                                                                                                                                                                                    ,        	                                                                                                                                                                                                           -                                                                                                                                                                                                                                 .          
                                                                                                                                                                                                   
             ,                                                                                                                                                                                                                              .           
                                                                                                                                                                                                        .                                                                                                                                                                                                                                    
     .                                                                                                                                                                                                                       	          .               
                                                                            	                                                                                                                                 -                                                                                                                                                                                                                  .                                                                                                                                                                                                                      1         .    	                                                                                                                                                                                                               -                                                                                                                                                                                                                   /                                   	                                                                                                                                                                                  0                                                                                                                                                                                                                     -                                                                                                                                                                                                                          -           	                                                                                                                                                                                                                  -                                     
                                                                                                                                                                                               0                                
                                                                                                                                                                                 /                               	                                                                                                                                                                                                    -                                                                                                                                                                                                                                     /                                                                                                                            
                                                                               1                                                                                        
                                                                                                                         ,                            
                                                                                                                                                                                                     .                                                                                                                                                                                                                1                                                                                        
                                                                                                                             0                                                                                       	                                                                                                                          0                                                                                                                                                                                                                     /                                                                                                                                                                                                    1                                                                                                                                                                                                       
0                                                                                                                                                                                                      1                                                                                                                                                                                                                -                                                                                                                                                                                                                                 0                                                                                                                                                                                              /                                                                                                                                                                                                                   -             
                                                                                                                                                                                                                ,                                                                                                                                                                                                                              -                                                                                                                                                                                                     	       -                                                                                                                                                                                                                     ,        	                    	                                                                                                                                                                                                      ,                                                                                                                                                                                                                            -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                    .                                                                                                                                                                                                                            ,                                                                                                                                                                                                               /                                                                                                                                                                                                             .                                                                                                                                                                                                                     .                                                                                                                                                                                                                        ,         
                                                                                                                                                                                                                     ,                                                                                                                                                                                                                          ,                                                                                                                                                                                                                
                     /                     	                                                                                                                                                                                                      ,                                                                                                                                                                                                               	                ,                
                                                                                                                                                                                                 .                                                                                                                                                                                                                 
                    .    
      
                                                                                                                                                                                                                   /                                                                                                                                                                                                                         -                                                                                                                                                                                                                        .                                                                                                                                                                                                                       +         -                          	                                                                                                                                                                                        .                                                                                                                                                                                                                  .                                                                                                                                                                                                              .                                                                                                                                                                                                               -                                                                                           	                                                                                                                                  -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                 /                                                                                                                                                                                                                 .               
                                                                                                                                                                                                            ,                                 	                                                                                                                                                                                                 0                                                                                                                                                                                                       
2                                                                                                                                                                                                               ,                               
                                                                                                                                                                                               2                                                                                                                                                                                                             1                                                                                  
                                                                                                                      0                          	                                                     	 	                                                                                                                               0                                                                                           	                                                                                                                          1                                                                                                                                                                                                                2                                                                                                                                                                                                     1                                                                                                                                                                                                     .                                                                                                                                                                                                               -                
                                                                                                                                                                                                                        2                                                                                                                                                                                                 	/                                                                                                                                                                                 
                            /                                                                                                                                                                                                                 -                                                                                                                                                                                                                           /                                                                                                                                                                                                                     /                                                                                                                                                                                                                 -           
                                                                                                                                                                                                                -                                                                                                                                                                                              	                          /                                                                                                                                                                                                                             -                                                                                          
                                                                                                                             /         
                                                                                                                                                                                                                         .                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                  ,                                                                                                                                                                                                     
                           -                                                                                                                                                                                                                   	             ,                                                                                                                                                                                                                    -             
                                                                                                                                                                                                     
                 .                                                                                                                                                                                                                      ,                                                                                                                                                                                                                       
               ,                                                                                                                                                                                                                                 -                
                                                                                                                                                                                                    
                   -                                                                                                                                                                                                                            -                                                                                                                                                                                                                                	     ,                                                                                                                                       	                                                       	                                  /                                                                                                                                                                                                                                  -                                  	                                                                                                                                                                                
                  -                                                                                                                                                                                                                              .                                                                                                                                                                                               	                         -                                                                                                                                                                                                                   	  -                                                                                                                                          	                                                                                         ,                                                                                                                                          
                                                                                           ,                                                                                                                                                                                                                 
               -                                                                                                                                                                                                                                     ,                                                                                                                                 	                                                                                  .                                                                                                                                                                                                                          -                                                                                                                                                                                                                                  -                                                                                                                                                                                                                                .                                 	                                                         
                                                                                                                                 -       	                                                                                                                                                                                                                          -                                                                                                                                                                                                                 	               -                                                                                                                                                                                                                                      ,                                      $                                                                                                                                                                                                     ,                                   
                                                                                                                                                                                                    .                                                                                                                                              	                                                                                
   ,                                                                                                                                                                                                        %                               ,                    
                                                                                                                             $                                                                                                    ,                     	                                                                                                                                                                                                               ,                                                                                                                                                                                                                        
             ,            	                                                                                                                          	                                                                                             .                                    	                                                                                                                                                                           	     
  ,                                                                                                                                                                                                                                            ,                                                                                                                                                                                                 	             
           
    
    ,                       	                                                                                                                                                                                                                  .                                                                                                                                	                                                                           	             -          	                                                                                                                                                                                                            .                                                                                                                                                                                                                          -       	      
                                                                                                                                                                                                                  -           	                                                                                                                                                                                                                    
    -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                    
                                 .                                                                                                                                                                                             	                                     ,        
                       	                                                                                                                                                                                  ,                                                                                                                                                                                                                       
           -           	                       
                                                                                                                                                                              
              -               	                                                                                                                                                                                                            
        -                                                                                                                                                                                                                        	-                                                                                                                                                                                                                         .                                   
                                                                                                                                                                                    -                                                                                                                                                                                                                         	                 0                                   	                                                                                                                                                                                         .                          	                                                                                                                                                                                                              
     ,                                                                                                                                                                                                                                           -                                                                                                                                                                                                                                  ,               
                                                                                                                                                                                                       	.                                                                                                                                                                                                                               	        ,                                                                                                                                                                                                                        .                                                                                                                                     	                                                                                       ,                                                                                                                                                                                                                                -                                                                                                                                                                                              
                                   -                                                                                                                                                                                                        
                                      -                                                                                                                                                                                                                                             -                                                                                                                                                                                                                        
     -                                                                                                                                                                                                                          ,                                    	                                                                                                                                                                          	                         ,                                       
                                                                                                 
                                                                                            
.                                                                                               	                                                                                                                          .                                                                                                                                                                                                                           -                                
                                                        	                                                                                                                              ,                                                                                                                                                                                                                              	,                                                                                                                                                                                                                                      ,                                                                                         
                                                                                                                                        
,                                                                                                                                                                                     	                               
.                                                                                                                                                                                                     
                            	-                                                                                                                                                                                                   	                                 -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                         

         	      ,                                                                                                                                                                                                                                  -                                                                                                                                                                                             	                                -            
                                                                                                                   	                                                                                        -                                                                                                                                                                                                                                       ,                
                     
                                                                                                                                                                             	                   /                                                                                                                                                                                                                         0                                                                                                                                                                                                                          ,                                                                                                                                                                                                                            #               -       	                                                                                                                                                                                                                            -                                                                                                                                                                                                                                 	    ,           
       	          	                                                                                                                                                                                                  ,                                                                                                                                                                                                            	                       
        -                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                            .                                                                                                                                                                                                                      
                  ,                                                                                                                                                                                                                                           ,                                                                                         
                                                                                                                     	              -                                                                                                                                                                                                                                         -                                                                                                                                                                                                                                  ,                                                                                                 
                                                                                                                              ,                                                                                                                                                                                                                                  	     .                                                                                                                                                                                                                               .                                                                                                                                                                                                                            ,                                                                                                                                                                                                                              

                .                                                                                                                                                                                                                             .                                                                                                                                                                                                                         -                                                                                                                                                                                                                              %    	      -                                                                                                                                                                                                                            
     ,                                      
                                                                                                                                                                                              -                                                                                                                                                                                                   
                             
        ,                                                                                                                                                                                                                                                   .                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                 .                                                                                                                                                                                                                -                                                                                                                                                                                                                               	     ,                                                                                                                                                                                                                                      	       ,                 0                                                                                                                                                                                                                          .                                                                                                                                                                                                                              .        
                                                                                                                                                                                                               ,                                                                                                                                                                                                                                            -         
                                                                                
                                                                                                                                            ,                                                                                              	                                                                                                                                        ,                                  $                                                                                                                                                                                                        ,                                                                                                     
                                                                                                                                    	,                                                                                                                                                                                                                                    ,            
                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                            .                                                                                                                                                                                               
                
          
    ,              	                                                                                                                                                                                                          -                                                                                                                                                                                                                 
            #      	    ,                                                                                               
                                                                                                                                           /                                                                                                                                                                                                                           -                       	                                                                                                                                                                                                       -                                                                                                                                                                                                                                   ,                                                                                                                                            
                                                                                         .                                                                                                                                                                                                                              ,                                 %                                                                                                                                                                                                -                                     	                                                                                                                                                                                                      -                                                                                                                                                                                                                                  -                                                                                                                                                                                                                                
.               
                                                                                                                                                                                                              ,                                                                                                                                                                                                                                  -                                                                                                                                                                                                                                          ,                                                                                                                                          
                                                                                      ,                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                            -                                                                                                                                                                                                                  
               -                                                                                                                                                                                                                            -                                                                                              	                                                                                                                                      ,            
                                                                                                                                                                                                                 -                                                                                                                                                                                                                     .                                                                                                                                                                                                                              .                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                           -                                                                                                                                                                                                      
                                  -                        	                                                                                                                                                                                                                   ,                                                                                                                                                                                                                          
                          -                                                                                                                                                                                                                                             -                                                                                                                                                                                                                 
     	    ,                
                                                                                                                                                                                 	                                    ,                                                                                                                                                                                                                                   ,                ,                                    	                                                                                                                                                                                                            -                                                                                                                                                                                                                                -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                            -                                                                                                                                                                                                                                        ,                                    #                                                                                                                                                                                                               ,                                         
                                                                                                                                                                                               ,                                                                                                                                                                                                                                                -                                                                                                                                                                                                                                         
,                                                                                                                                               ,                                                             
                                       -                                                                                                                                                                                          	                                ,                                                                                                                                                                                                                                   "          ,           )                                                                                                                                                                                                                                 -                                                                                                                                                                                              
                        
     ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                 -                                      
                                                                                                                                                                                             .                                                                                                                                                                                                            	          	  .                     
                                                                                                                                                                                           
               -                                                                                                                                                                                                                                  ,                 	                                                                                                                                                                                                                           ,                                                                                              	                                                                                                                               	     -                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                         ,                                                                                                                                                                                             
                                  -                                                                                                                                                                                                                     	       /           	                                                                                                                                                                                                      
               ,                                                                                                                                                                                                                         -                                                                                                                                                                                                                               ,                                                                                                                                                                                                              
.                                                                                                                                                                                                                          -        	                                                                                                                                                                                                                 ,                                                                                                                                                                                                                              -                               	                                                                                                                                                                                        .                                                                                                                                                                                                                                   
   -                                                                                                                                                                                                                  -                                                                                                                                                                                                              	                 ,                                                                                                                                                                                                                                .                                                                                                                                                                                                                               -                                                                                                                                                                                                                      	           ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                          	                              -                    	                                                                                                                                                                                               -                                                                                                                                                                                                                       
    ,                 $       	                                                                                                                                                                                                              -                                                                                                                                                                                                                           
   -                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                   )              ,         	      	       
                                                                                                                                                                                                        -                                                                                                                                                                                                                	    -                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                         ,                                                                                                
                                                                                                                                             -                                          	                                                                                                                                                                                               -                                      %   
                                                                                                                                                                                             ,                                                                                                                                                                                                                            
           ,                     	                                                                                                                                                                                      	                                     ,                                                                                                                                            	                                                                                         -                                                                                                                                                                                                                             ,                                                                                                                                                                                                                             .     	   ,                                                                                                                                                                                                                                       ,           
                                                                                                                                                                                                              -                                                                                        
                                   	                                                                                             /                                                                                                                                                                                                                         	    ,          %                                                                                                                                                                                                                              -                                                                                                                                                                                                                       -                                                                                                                                    
                                                                                             	-                                                                                                                                                                                                                       	         ,                                                                                                                                                                                                                                       .                                                                                                                                                                                                                                -      
  
                                                                                                                                                                                                               ,                                                                                                                                                                                                                           	      ,                                  	                                                                                                                                                                                         -                                                                                                                                                                                                                  .                                                                                                                                                                                                          
                -                                                                                                                                                                                                                  -                                                                                                                                                                                                                                    -                                                                                                                                                                                                                          -                                                                                                                                                                                                                               -                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                            /         	                                                                                                                                                                                                         .                                                                                                                                                                                                                                  -                                                                                                                                                                                                                           -              	                                                                                                                                                                                                        	            .                                                                                                                                                                                                        	           .          
                                                                                                                                                                                                                        ,                                                                                                                                                                                            	                           /                 
                                                                                                                                                                                                                 -                                                                                                                                                                                                 	                                    -                                                                                                                                                                                                                                     -                                                                                                                                                                                                                                ,      	             &                                                                                                                                                                                                                             -                                                                                                                                                                                                                        -                                                                                                                                                                                                                                    /                                                                                                                                                                                                                 	                      ,                  	                                                                                                                                                                                                                    	.                                                                                                                                                                                                                         .                	                                                                                                                                                                                                        -                                                                                                  
                                                                                                                                          -                                                                                                                                                                                                                                            	-                                     0                                                                                                                                                                                                      ,                                  	                                                    	                                                                                                                                          ,                                                                                                                                                                                                       # 	                             ,                                                                                                                                                                                                          !                                   ,                                                                                                                                          $                                                                                                ,                                     
                                                                                                                                                                                              ,                                                                                                                                                                                                                            	
              ,                                                                                                                                                                                                                                   -                                                                                                                                                                                                                
       -                                                                                                                                                                                                                               .                                                                                                                                                                                                                               
      ,             2                                                                                                                                                                                                                             .                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                       .                                                                                                                                                                                                                           ,                                                                                                                                 	                                                                                                -                                                                                            	                                                                                                                                          -                                                                                                                                                                                                                                   /                                                                                                                                                                                        	                              ,                                                                                                                                                                                              	                                     ,                                                                                                                                                                                                                                 	 -                   
                                                                                                                                                                                                      /                                                                                                                                                                                                               .       	   
                                                                                                                                                                                                             -                                                                                                 
                                                                                                                                     2                                                                                                                                                                                                            .                                                                                                                                                                                                               .                                                                                                                                                                                                                                      ,                                                                                                                                                                                                                         	  1                                                                                                                                                                                                           0                                                                                                                                                                                                         .                                                                                                                                                                                                                               ,                                                                                                                                                                                                                          /                                                                                                                                                                                                                           ,                                                                                                                                                                                                                       -                                                                                                                                                                                                                                      .                                                                                                                                                                                                     	         -                                                                                                                                                                                                                      .                                                                                                                                                                                                                         
         ,                                                                                                                                                                                                                .                                                                                                                                                                                                           -    
                                                                                                                                                                                                                   /                                                                                                                                                                                                                         ,             	'                                                                                                                         
                                                                                               -                                                                                                                                                                                                               ,                                                                                                                                                                                                                       .                                                                                         
                                                                                                                          /                                                                                                                                                                                                                                -                                  	                                                                                                                                                                                       .                                                                                                                                                                                                                          2                                                                                                                                                                                                      /                                                                                                                                                                                                                    	    ,                                                                                                                              	                                                                                     .                                                                                                                                                                                                                    .                                                                                                                                                                                                                      "      /                                                                                                                                                                                                                            /                                                                                                                                                                                                            -                                                                                     
                                                                                                                                   .                                                                                                                                                                                                          
      -                                                                                                                                                                                                                  1                                                                                                                                                                                                                .                                                                                                                                                                                                                               .                                                                                                                                                                                                                .                                                                                                                                                                                                                 .                                                                                                                                                                                                                                -        	                                                                                                                                	                                                                                        -                                                                                                                                                                                                       .                                                                                                                                                                                                            -                                                                                                                                                                                                                
                 .                                                                                                                                                                                                        	2                                                                                                                                                                                                     -                                                                                                                                                                                                                                -                                                                                                                                                                                                                  
   .                                                                                                                                                                                                           .                               	                                                                                                                                                                             -                                                                                                                                                                                                                           0                                                                                                                                                                                                        /                                                                                                                                                                                                         	        1                                                                                                                            	                                                     	                            /                                                                                                                                                                                                  	         /                                                                                                                                                                                                                 	/      
                                                                                                                                                                                                                .                                                      	                                                                                                                                                              .                                     
                                                                                                                                                                                               .                                                                                                                                                                                                                        -   	                                                                                                                                                                                                                            /                                                                                                                                                                                                                      ,                                                                                                                                                                                                                     	     /                                                                                                                      
                                                                                       .             
                                                                                                                                                                                                                   -                                                                                                                                                                                                                                        ,                
                                                                                                                                                                                                              /                                                                                                                                                                                                                        ,                              	                                                                                                                                                                                                -                                                                                                                                                                                                                               -             
                                                                                                                                                                                                               0                                                                                                                       	                                                                                      .                                                                                                                                                                                                                .                                                                                                                                                                                                         	,                                                                                        
                                                                                              	                       
      .                                                                                                                                                                                                                  -                                                                                                                                                                                   
                              -                                                                                                                                                                                                                         
   -                               	                                                                                                                                                                                    0                                                                                                                                                                                                               -                                                                                                                                                                                                                        /                                                                                                                                                                                                                                   .                                                                                                                                                                                                  
                 1                                                                                                                                                                                                                   /                                                                                                                                                                                                                                   /                       
                                                                                                                                                                                              
                /                                                                                                                                                                                                                      -                                                                                                                                                                                                                                   -             	                                                                                                                                                                                                                   /                                                                                                                                                                                                                              0                                                                                                                                                                                                             1                                                                                                                                                                                                                        	    .                                                                                                                                                                                                                     0                                                                                                                                                                                                             -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                      /                                                                                                                                                                                                              -                                                                                                                                                                                                                      -                                                                                                                                                                                                                            .                                                                                                                                                                                                                	                 /                                                                                                                                                                                                              	              	   /                                                                                                                                                                                                     0  
   
                                                                                                                                                                                                                  -                                                                                                                                                                                                                                   0                                                                                                                                                                                                                    /                                                                                                                                                                                                          /                                 	                                                    	                                                                                                                              .                                                                                                                                                                                                                 -                                                                                                                                                                                                                          .                                                                                                                                                                                                                           .                                                                                                                                                                                                                /                                                                                                                           	                                                                             -                                                                                                                                                                                                                                 .                                                                                                                                                                                                                          .                                                                                                                                                                                                                        -                          	                                                                                                                                                                                     /   	     	                                       	                                                                                                                                                                              ,                                                                                                                                                                                                                                    .                                                                                                                                                                                                                            .                                                                                                                                                                                                                      2                                    	                                                                                                                                                                           0                                                                                                                                                                                                              1                                                                                                                                                                                  	                       -                                                                                                                                                                                                                          -                                                                                                                              	                                                                                      -                                                                                                                                                                                        	                           .                                                                                                                                                                                                                 .                                                                                                                                                                                                                 .                                                                                                                                                                                                                        /                                                                                                                                                                                                                          /                                                                                                                                                                                                                 .                                                                                                                                                                                                         ,                                                                                                                                                                                                                        -                                                                                                                                                                                                                    -                                                                                                                                                                                                                     -  	  	                                                                                                                                                                                                                     .      	                                                                                                                                                                                                                   -                                                                                                                                                                                                  &                              -                                                                                                                                                                                                                               -                                                                                                                                                                                                                                   -                                                                                                                                                                                                                            0                                                                                                                                                                                                                     .        
                                                                                                                                                                                                                  .                                                                                                                                                                                                                  /                                                                                                                                                                                                             2                                                                                                                                                                                                    -                                                                                                                                                                                                                       1                                                                                                                                                                                                        /                                                                                                                                                                                                                  /                                                                                                                                                                                                                     .     
                                                                                                                                                                                                              .                                                                                                                                                                                                     -                                                                                                                                                                                                                                  /                                  	                                                                                                                                                                                       0                                                                                                                                                                                                                                 /                                                                                                                                                                                                          
       ,           
                                                                                                                                                                                                                    .                                                                                                                                                                                                                         /                                                                                                                                                                                                              -                                                                                                                                                                                                      
          -                  
                                                                                                                                                                                                          .                                                                                                                                                                                                                    
   -                        
                                                                                                            
                                                                                              .                                                                                                                                                                                                                          .                                                                                                                                                                                                                              1                                                                                                                                                                                                                   0                                                                                                                                                                                                           /                                                                                                                                                                                                              /                                                                                                                                                                                                                        /                                                                                                                                                                                                           	0                                                                                                                                                                                                         .                                                                                                                                                                                                             
.                                                                                                                                                                                                             -                                                                                                                                                                                                                                
  /                                                                                                                                                                                                                  -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                         0                                                                                                                                                                                      	                    .                                                                                                                                                                                                         /                                                                                                                                                                                                
            	     -      
                                                                                                                                                                                                                            /                                                                                                                                                                                                                      	        0                                                                                                                                                                                                           ,                                                                                                                                                                                                                              0                                                                                                                                                                                                               /                                                                                                                                                                                           !                            	      /                 
                                                                                                                                                                                                         .                                                                                                                                                                                                           
        
    .                                                                                                                                                                                                                          .                                                                                                                                                                                                                              -                                                                                                                                                                                                              	                 .                                                                                                                                                                                                               .                                                                                                                                                                                                                    0                                                                                                                                                                                                        	-                                                                                                                                                                                                             	               0                                                                                                                                                                                                    
.                                                                                                                                                                                                                     .                                                                                                                                                                                                             	              -                                                                                                                                                                                                                        -                                                                                                                                                                                                          	   -           	                                                                                                                                                                                                                     .                                                                                                                                                                                                                     1                                                                                                                                                                                                              	               -                                                                                                                                     
	                                                                           
           ,            
                                                                                                                                                                                                        /              	                                                                                                                                                                                                            ,                                                                                                                                                                                                             
               /                                                                                                                                                                                                       
              -    
                                                                                                                                                                                                                          1                                                                                                                                                                                                                   ,                                                                                                                                                                                                                             .                                                                                                                                                                                                                              .                                                                                                                                                                                                                   -                                                                                                                                                                                                                        /                                                                                                                                                                                                            0                                                                                                                                                                                                          -                                                                                                                                                                                     	                                0                                                                                                                                                                                                             0                                                                                                                                                                                                   .                               	                                                                                                                                                                                    .                                                                                                                                                                                                                -                                                                                                                                                                                	                                          	   0                                                                                                                                                                                                               0                                                                                                                                                                                                                        -                                                                                                                                                                                                                                  /                                                                                                                                                                                                                       -                                                                                   	                                                                                                                              /                                                                                                                                                                                                                  -       	              	                                                                                                                                                                                                                   /                                                                                                                                                                                                         	              /                                                                                                                                                                                                              -      	                                                                                                                                                                                                                  .                                                                                                                                                                                                                            0                                                                                                                                                                                                                          /                                                                                                                                                                                                                   /                                                                                                                                                                                                                     #       .                                                                                                                                                                                                                  1                                                                                                                                                                                                                       -        	                                                                                                                                                                                                           /                                                                                                                                                                                                                          .               
                                                                                                                                                                                                              /                                                                                                                                                                                                            -         
                                                                                                                                                                                                    /                                                                                                                                                                                                             
            .                                                                                                                                                                                                                   
      
  /                                                                                                                                                                                                        	.       	                                                                                                                                                                                                          .                                                                                                                                                                                                                &           .            	                                                                                                                                                                                                      -                                                                                                                                                                                                                     -                                                                                                                                                                                                                           .                                                                                                                                                                                                              /             	                                                                                                                                                                                                                 /                                                                                                                                                                                                                      	   /                                                                                                                                                                                                                	/                                                                                                                                                                                                     
          ,     
                                                                                                                                                                                                                                /                                                                                                                                                                                                              	       ,                                                                                                                                                                                                                                -                                                                                                                                                                                                                %               ,                                                                                                                                                                                                                            .                                                                                                                                                                                                                1                                                                                                                                                                                                            /                                    
                                                
                                                                                                                            -                                                                                                                                                                                                                         1                                                                                                                                                                                                      0                                                                                                                                                                                                    -                                                                                                                                                                                                               .                                                                                                                                                                                                         
,                                                                                                                                                                                                                             .  
           
       
                                                                                                                                                                                               0                                                                                                                                                                                        
                              ,                                                                                                                                                                                                                                            1                                                                                                                                                                                                                  /                                                                                                                                                                                                               .                                                                                                                                                                                                         
         ,          ,                                                                                                                                                                                                                                 .                                                                                                                                                                                                          
           /                                                                                                                                                                                                             -                                                                                                                                                                                                                 -                                                                                                                                                           	                                                           -                                                                                                                                                                                                                              .     	                                                                                                                                                                                                             /                                                                                                                                                                                                                      /            
                                                                                                               	                                                                                       ,                                                                                                 "                                                                                                                                                .                                                                                         
                                                                                                                                   ,                                                                                                                                                                                                                 	       *              0                                                                                                                                                                                                                              -                                                                                                                                                                                                              -                                                                                                                                                                                                                            	  
     -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                  	         	   ,                                                                                            
                                     
                                                                                          .                                                                                                                                                                                                         1                                                                                                                                                                                                                       .                          	                                                                                                                                                                                       ,                                                                                                                                                                                                            
       /                                                                                                                                                                                                                .                                                                                                                                                                                                                       /                                                                                                                                                                                                                    -                                                                                                                                                                                                   
                
  -                                                                                                                                                                                                                         /                                                                                                                                                                                                            1                                                                                                                                                                                                                    -                                                                                                                                                                                                                     .             ,      
            '                                                                                                                                                                                                                       1                                	                                                                                                                                                                           ,                                                                                                                                                                                                           2                                                                                                                                                                                                                -                                                                                               '                                                                                                                                         -                        
                                                                                                                                                                                         .                               
                                                                                                                                                                                              3                                                                                                                                                                                                           	.                                                                                                                                                                                                                       0                                                                                                                                                                                                           0                                                                                                                                      	                                                         
                            0                                                                                                                                                                                                                   -              	                                                                                                                                                                                                                     0                                                                                                                                                                                                            .                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                    /                                                                                                                                                                                                     1                                                                                                                                                                                                               /                                                                                                                                                                                                                    	               .                                                                                                                                                                                                                   -                                                                                                                                                                                                           	                    /       	   
                     	                                                                                                                                                                                     .                                                                                                                                                                                  
                                    /                                                                                                                                                                                                    .                                                                                                                                                                                                                        2                                                                                                                                                                                                       .                               	                                                                                                                                                                                       -        	     
                                                                                                                                                                                                              -                                                                                                                                                                                                                	         	        .                                                                                                                                                                                                                           	      2                                                                                                                                                                                                                 .                                                                                                                                                                                                                            ,                                                                                                                                                                                                                
                    ,                                                                                                                                                                                                         
                 
    /                                                                                     	                                                                                                                            1                                                                                                                                                                                                    	.                                                                                                                                                                                                                      .                                                                                                                                                                                                              .                                                                                                                                                                                                                   	      .                                                                                                                                                                                                                             ,                                                                                                                                                                                                                  /              	                                                                                                                                                                                                             -                                                                                                                                                                                                                            -              %                                                                                                                                                                                                             -                                                                                                                                                                                                             .   	           
                                                                                                                                                                                                                 -                                                                                                                                                                                                                        ,                        	                                                                                                                                                                                                            0                                                                                                                                                                                                                 -                                                                                                                                                                                                              .                                                                                     	                                                                                                                    .                                                                                                                                                                                                                                  /                                                                                                                                                                                                                           1                                                                                                                                                                                                                              1                                                                                                                                                                                                 	-                                                                                                                                                                                          
                                /                                                                                                                                                                                      	 
                               /                                                                                                                                                                                                                      .                                                                                                                                                                                                                         -                                                                                                                                                                                                                                       0                                                                                                                                                                                                                          -                                                                                                                                	                                                                                           -                                                                                                                                                                                                                                  ,                                        	                                                                                                                                                                                            /                                                                                                                                                                                                                   0   	            
                                                                                                                                                                                                              -                                                                                                                                                                                                                                     -                                                                                                                                                                                                             -                                                                                                                                                                                                                          ,                                	                                                                                                                                                                                            .                                                                                                                                                                                                                 /                                                                                                                                                                                              -                                                                                                                                                                                                                              
  /                                                                                                                                                                                                                   ,                              
                                                        
                                                                                                                                  ,         	                                                                                                                                                                                                                    /                                                                                                                                                                                                                         #	            	    -                                                                                                                                                                                                                                 0                                                                                                                                                                                                             ,                                                                                                                                                                                                                                  /                                                                                                                                                                                                               	                   -                                                                                                                                                                                                                             	  .                                                                                                                                                                                                                       .                                                                                                                                                                                                          .                                                                                                                                                                                                                        
       -      	  	                                                                                                                                                                                                                -                                                                                                                                                                                  	                              -                                                                                                                                                                                                                      -                                                                                                                                                                                                                     -          
                                                                                                                                                                                                    /                                                                                                                                                                                                  
                     ,                                                                                                                                                                                                                             .                                                                                                                          	                                                                                         -                   	                                                                                                                                                                                                     /                                                                                                                                                                                                             $             -                      	                                                                                                                                                                                                         /                               	                                                                                                                                                                                     1                                                                                                                                                                                                              /                                                                                        
                                                                                                                      .                                                                                                                                                                                                                                      .                                                                                                                                                                                                                          .                                  
                                                                                                                                                                                               2                                                                                                                                                                                                             .                                                                                                                                     
                                                    	                        .                                                                                                                                                                                                                            -                                                                                               	                                                                                            
                             /                                                                                                                                                                                                                 ,                     
                                                                                                                                                                       	                                      0                                                                                                                                                               	                   
                                /            
                                                                                                                                                                                                         .                                                                                                                                                                                                                          
     "       ,         !                                                                                                                                                                                                                               .                                                                                                                                                                                                              /    
 	                                                                                                                                                                                                                  .                                                                                                                                                                                                                       
       0                                                                                                                                                                                                                 .    
                                                                                                                                                                                                                      -                                                                                                                                                                                                                      /                                                                                                                                                                                                                                 
        ,             	                                                                                                                                                                                  
                                 ,                                    
                                                                                                                                                                                       -                                                                                                                                                                                                    	                         
      	      ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                      -                                                                                                                                                                                                                                  -                                                                                                                                                                                                                            .                                                                                                                                                                                                                              .                                                                                                                                                                                                                               -       
                          	   	                                                                                                                                                                                      .                                                                                                                                                                                                                                 	    ,                                                                                                    	                                                                                                                      !                ,          	                                                                                                                                                                                                                                 ,                                                                                                                                                                                                                         	          -                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                       
        -                   
                                                                                                                     !                                                          	                                     ,                                                                                                                                                                                                                                  	   -                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                              ,                                                                                                                                                                                                       	                                 .                                                                                                                                                                                                                              .                                                                                                                                                                                                                      ,                                                                                                                                                                                                                           
    -        	                                                                                                                                                                                                                      -                	                                                                                                                                                                                                        /           
                     
  	                                                                                                                                                      	                                  ,                                                                                                                                                                                                                                       ,                                   !                                                                                                                                                                                           .                 	                                                                                                                                                                                                                    -           
                                                                                                                                                                                                                       ,                                                                                                                                                                                                                      	            ,                                                                                                                                                                                                                                  .                                                                                                                                                                                         
                    
         0                                                                                                                                
                                                                                     ,                                                                                                                                                                                                                            !    
      -                                                                                                                                                                                                                                .                                                                                                                                                                                                                            /                                                                                                                           	                                                                                          ,                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                 .                                                                                                                                                                                                                           	.        
                                                                                                                                                                                                             ,          	                                                                                                                                                                                                                                  -                                                                                                                                                                                                                                   .                                                                                                                                                                                                                                    ,                                                                                       
                                                                                                                                   -                                                                                                                                                                                                  
                                 -                                                                                                                                    
                                                                                        ,                                                                                                                                                                                                                              -                                                                                                                                                                                                                     	         -                                                                                                                                                                                                                        ,       .                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                  
         !         -            
     
                                                                                                                                                                                                           	        ,                                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                   ,                                                                                                                                                                                                                                          .                                                                                                                                                                                                                                       -                                                                                                                                                                                                                           -                                                                                                                                                                                                                            ,                                                                                                                                                                                                                          -                                                                                                                                                                                                                    	    
     -                                                                                                                                                                                                                           .                                                                                                                                                                                                                           .                                                                                                                                                                                                                            
     -                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                               ,                                                                                                                                          	                                                                                             0                                                                                                                                                                                                                     -                                                                                                                                                                                                                         ,                                                                                                                                                                                                                             $             ,           
                                                                                                                             

                                                                                                ,                                                                                                  	                                                                                                                                     -          $                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                              
         
      	  ,                                                                                                 & 	                                                                                                                         	                  ,                                 )                                                                                                                                                                                                         ,                                      )                                                                                                                                                                                                  ,                                                                                                                                                                                                           	                                 
     ,                                                                                            
                                                                                                                                       ,            	                                                                                                                                 $                                                                                         ,                                                                                                                                               1                                                                                                  -                                                                                                                                                                                                                       
                        ,             (              	                                                                                                                                                                                                                       -                                                                                                                                                                                                                 	              ,                       	                                                                                                                                                                                                         .                                                                                                
#                                                                                                                                          ,                       
                                                                                                                                                                                               	              -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                         .                                                                                                                                       &                                                                                            -                                                                                                                                                                                                                                 -                                                                                                                                                                                                                            .                                                                                                                                                                                                                                         -      
                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                    -                                   	                                                                                                                                                                            .                                                                                                                                                                                        	                                        ,                                                                                                                                                                                                                                 -                                                                                                                                                                                                                                    ,                                                                                                                                                
                                                                                          .                                                                                                                             	                                                                                             ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                       /                                                                                                                             	                                                                                            .                                                                                                                                                                                                                          ,                                 	                                                                                                                                                                                                   ,                                                                                                                                                                                                   
                                 /                                                                                                                                                                                                                            ,                                   1                                                        	                                                                                                                                         .                                                                                                                                                                                                                                     .                                                                                                                                                                                                             -                                                                                                                                                                                                                            ,                                                                                                                                                                                                                                        -        -                	                                                                                                                                                                                                          -                                                                                                                                                                                                                	             /                                                                                                                                                                                                                      ,                                                                                                                                                                                                                                )                -                                                                                                                                                                                                                         ,                                                                                                                                                                                                              
               
                 -                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                  "             
     ,                                                                                                      &                                                                                                                                            .                                                                                                                                                                                                                           .                                                                                                                                                                                                                                ,                                                                                                                                                                                                              
                     
                 ,                                                                                                                                                                                                                                              "         -                                                                                                                                                                                                                            /                                                                                                                                                                                                                         ,                                                                                                                                                                                                                                        
     .                                                                                                                                                                                                                            ,                                                                                                    	                                                                                                              
               ,              	                                                                                                                                                                                                             ,                                                                                                                                                                                                                               .                                                                                                                                                                                                                         -                                                                                                                                                                                                                                      -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                                       .             	                                                                                                                                                                                                
             -                                                                                                                                                                                                                      .             
                                                                                                                                                                                                      ,                                                                                                                                                                                                                            -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                      	   ,           	                                                                                                                                                                                                          	                ,                                                                                                                                                                                                                                           -                                                                                   	                                                                                                                    	              ,                                                                                                                                                                                                                                 -                                      	                                                                                                                                                                                             ,                                                                                                                                                                                                                                                .                                                                                                                                                                                                                                .                                                                                        
                                                                                                                                   -                                                                                                                                                                                                                       -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                             /                                                                                                                                                                                                                          .                                                                                                                                                                                                                            ,                                                                                                                                                                                                        
              ,           "    	                                                                                                                                                                                                                     -                                                                                                                                                                                                                      -            
                                                                                                                                                                                                                        ,                                                                                                                                                                                                                                      	   	
   -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                     
  -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                               -              #                                                                                                                     
                                                                                        .                                                                                                                                                                                                              ,                                                                                                                                                                                                                                ,                                                                                                   
                                                                                                                             
    ,                                                                                         	                                                                                                                                    -                                                                                                                                                                                                                  .                                -                                                                                                                                                                                               ,                                                                                                                                                                                                                                         ,                                                                                                       
                                                                                                                                    ,                                                                                                                                                                                                                             ,                                   %                                                                                                                                                                                                       -                                                                                                                                                                                                                                           -          
                                                                                                                                                                                                        	           	    -                                                                                             	                                                                                               
                                   -                                                                                                                                                                                                                                    ,                                                                                                                                                                                                                             
              -                                                                                                                                                                                                                                       /                                                                                                                                                                                                                           ,                                                                                                                                                                                                                	                    ,                                                                                                                                                                                                               ,                                                                                            	                                                                                                                                          -                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                  ,                                                                                                                                                                                                   $                                   ,                 	                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                                .                                                                                                                                                                                                                               1            ,                                                                                                                                                                                                                                   	   	     ,                    	                                                                                                                                                                                                                  ,                                                                                                                                                                                                                           
             .                                                                                                                                                                                                                                 
      ,                                                                                                                                                                                                                   	            -                                                                                                                                                                                                                             %             ,             (       
                                                                                                                                                                                                               	          ,                        	                                                                                                                                                                                                         "        -                                                                                                                                                                                                                             ,      	                                                                                                                                                                                                                                   ,               )                                                                                                                                                                                                                          .                                                                                                                                                                                                                      -                  /                                                                                                                                                                                                                   ,                                                                                         	                                                                                                                                    ,             
                          4                                                                                                                                                                                                            ,                                      2                                                                                                                                                                                                                ,                                    >                                                                                                                                                                                                  ,                                                                                                                                                                                                                                             -                                                                                                                                                                                                                                   ,                                                                                                                                       
                                                                                                ,                                             
                                                                                                                                                                                                        -            !                                                                                                                                                                                                                       0                                                                                                                                                                                                            	        -             	                                                                                                                                                                                                                ,                                                                                                                                                                                                                                    ,       	                                                                                      (                                                                                                                                                   ,                                                                                              
                                                                                                                                       ,                                 +                                                                                                                                                                                                      ,                        
                                                                                                                                                                             
                                        ,                                                                                                                                                                                                                                            	 ,                                         	                                                                                                                                                                                                    ,                                                                                                                                                .                                                                                              ,                                                                                                                                             '                                                                                           ,           
                                                                                                                                                                                                                               -                                                                                                                                                                                                 	                             -                                                                                                                                                                                                                -                                                                                                                                                                                                
                                -                                                                                                                                                                                                                         .                                                                                                                                                                                                                    -                                                                                                                                                                                                                        /                                                                                                                                                                                                                       ,                                                                                         
                                                                                                                                     ,      
                                                                                                                                	                                                                                                    ,          	                                        	                                                                                                                                                                                       .                                                                                                                                                                                                      %                                      ,                                                                                                                                                                                                                         ,                                                                                                                                                                                                                             
/                                                                                                                                                                                                                                          ,                                                                                                                                                                                                                                     /                                                                                                                                                                                                                                  ,                                                                                                                                                                                                                             	/                                                                                                                                                                                                                                        ,                                                                                                                                                                                                   
                                ,                                                                                                                                                                                                                                !           -                                          	                                                                                                                                                                                   	           -                                                                                                                                                                                                                            
    ,                                                                                                                                                                                                                                         ,             	                        	                                                                                                                                                                                          ,                                                                                                                                                                                                                                              
 .                  
                                                                                                                                                                                                                                -                                                                                                                                                                                                                          ,         
                                                                                                                                                                                                                                      -                                                                                                                                                                                                   
                              	   ,                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                             ,                8                                                                                                                                                                                                                           -                                                                                                                                                                                                                                   
      -                                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                   	                  ,                                                                                                                                                                                                                      ,         
                                                                                                                                                                                                                    ,                                                                                                                                                                                                                                               -                                    1                                                                                                                                                                                                       ,                                          =                                                                                                                                                                                                               ,                                      B                                                                                                                                                                                                                 ,                                                                                                                                                                                                                                  ,                                                                                                                                     	                                                                                      ,                                                                                                                                                  >                                                                                                     ,                                                                                                                                                                                                                                           
,                                                                                                                                                                                                                               ,                                                                                                                                                                                             
                          
       ,                                                                                                                                                                                               
                                  ,                                                                                                                                                                                                                                            ,               	                 
                                                                                                                                                                                                ,                                                                                                                                                                                                                                  .                                                                                                                                                                                                                                       ,        
                                                                                                                                                                                                                                        ,                                                                                                                                                                                                                               ,             	      &                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                             ,                                                                                                                                                                                                                                                  -                                  
                                                                                                                                                                                           -                                                                                                                                                                                                                            0                                                                                                                                                                                                                 -         	     
                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                      -                                                                                                                                                                                                                           ,             
                                                                                                                                                                                                         -          	                                                                                                                                                                                                                               -                                                                                                                                                                                                                                     -           
    	                                                                                                                                                                                                              ,                                                                                                                                                                                                                            .                                                                                                                                                                                                                                "           .             
                                                                                                                                                                                                                 ,                                                                                                                                                                                                                 -                                                                                                                                                                                                                 -                 
                                                                                                                                                                                                                           ,                                                                                                                                	                                                                                            ,                                                                                                                                                                                                                     	         .                                                                                                                                                                                                                            , 
                	                                                                                                                                                                                                             /                                                                                       
                                                                                                                                 /     	                
                                                                                                                                                                                                                 .                                                                                                                                                                                              	                            	    ,                                                                                                                                                                                                                          ,                                     
                                                                                                                                                                                               /                                                                                                                                                                                                                            .                                                                                                                                                                                                              	         	    /                                                                                                                                                                                                            ,        
      
       	                                                                                                                                                                                                           -                                                                                                                                                                                                                                   .                                                                                               
                                                                                                                               /                                                                                                                                                                                                                           -        	   	                                                                                      
                                                                                                                                       -                                                                                                                                                                                                                            -                                                                                                                                                                                                                                 ,                                   	                                                                                                                                                                                        -                                                                                                                                                                                                                          .                                     	                                                                                                                                                                                                    .                                                                                                                                                                                                                          -           
                                                                                                              
                                                                                         ,                                                                                                                                                                                                                          ,                 	       	                                                                                                                                                                                                            -                                                                                                                                                                                                            ,                                                                                                                                                                                                                  	          ,               	                                                                                                                    
                                                                                                  -                                                                                                                                                                                                                      .                                                                                                                                                                                                                          -       
                         
                                                                                                                                                                                                     .                                                                                                                                                                                                                           
   /                                                                                                                                   	                                                                                         -                                                                                                                                                                                                                 -                                                                                                                                                                                                                                     ,                                                                                                                                                                                                                                         -                                                                                                                                                                                                                    *                     ,                                       
                                                                                                                                                                      	              .                                                                                                                                                                                                                        "      
             ,                                                                                                                                                                                                	                           .                                                                                                                                                                                                                                       ,                 	       	                                                                                                                                                                                      	                 .                                                                                                                                                                                                                
                            ,                                                                                                                                                                                                                                  ,           	             	                                                                                                                                                                                                            .                                                                                                                                                                                                       	           -                                                                                                                                                                                                                        %                  ,                                                                                                                                                                                                                            ,         	                                                                                                                                                                                                                     .                                                                                                                                                                                                                 -                                                                                                                            
                                                                                               .                                                                                                                                                                                                                ,            !                                                                                                                                                                                                                                      /           
                                                                                                                                                                                                                 -        
    	                                                                                                                                                                                                           -                                                                                                                                                                                                                          
                 ,                                                                                                                                                                                                                                           /                                                                                                                                                                                                                      ,        
                                                                                                                                                                                                               ,                                      
                                                                                                                                                                                                 ,                                                                                                                                                                                                                                    .                                                                                      	                                                                                                                        ,	                                                                                                                                                                                     	                                  ,                                                                                                                                                                                                               	              ,                                                                                                                                                                                                 
                                  -                                                                                                                                                                                                                     ,                                                                                                                                                                                                                          ,                                                                                                                                                                                                  	                           -        !                                                                                                                                                                                                                    1         	                                                                                                                                                                                
                                ,                                                                                                                                     
                                                                                         ,                                                                                                                                                                                                                                      .       !            	                                                                                                                                                                                                               0           
                                                                                                                                                                                                            -              	                                                                                                                                                                                                                        .                             	                                                                                                                                                                                     	,                                                                                                                                                                                                                                  -                                                                                                                                                                                                                        ,        	                                                                                                                                                                                                                  ,                                                                                                                                                                                                                                ,                                                                                                                                                                                                                           ,                                                                                                                                        	                                                                                .                                                                                                                                                                                                                              ,                                                                                                                                                                                                                     	            ,                                                                                                                                                                                                                                    -                                                                                                                                                                                                                ,                                                                                                                                                                                                                ,                                                                                                                                                                                                           	                         
     ,                   	                                                                                                                                                                                                    
                 .                                                                                                                                                                                                                    0                                                                                                                                                                                                         		    	         ,                                                                                                                                   		                                                                                       ,                                                                                           
                                                                                                                                   -                                                                                                                                                                                                                 	             .                                                                                                                                                                                                                       -                                                                                                                                                                                                                                       -          
                                                                                                                                                                                                                  ,           	                                                                                                                                                                                         
                                  ,                  $                                                                                                                        	                                                                                               ,                                                                                                                                                                                                                                     G             
       .                 *                                                                                                                                                                                                               /                                                                                                                          	                                                                             
          -                                                                                                                                                                                                                                     	,                                                                                                                                                                                                                             
       .                    .                                                                                                                                                                                                                               .                                                                                                                                                                                                                     ,                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                    
         ,                                                                                                                                                                                                                                     .          	                                                                                                                                                                                                                   0                                     -                                                                                                                                                                                                 ,                                                                                                                                                                                                                                               ,                                                                                                                                                                                                                            ,                                                                                                                                                                                                                              .                                                                                                                                           7                                                                                                    ,                                                                                                                                                                                                                                           3         /                                                                                                                                                                                                                      ,                                                                                                                                     
                                                                                   
    ,                                                                                                                                  	                                                                                            ,                                                                                                                                                                                                                                            ?            .            &                                                                                                                                                                                                                        /                                                                                                                                                                                                                ,                   
                                                                                                                                                                                                                  .                                                                                                                                                                                                                              .                                                                                                                                           	                                                                                         .                                                                                                                                                                                                                            ,                                                                                                                                                                                                                           -                              	                                                                                                                                                                                          -                                                                                                                                                                                                                          ,                                                                                                                                                                                                                
 .                     
                                                                                                                                                                                                                  ,                                                                                                                                                                                                    	                           -             
                                                                                                                                                                                               	                 /                                                                                                                           	                                                                                        .                                                                                                                                                                                                                                    ,                                                                                                                                                                                                	                            -              	                                                                                                                                                                                                                   
          ,              	                                                                                                                 
                                                                                             -                                                                                                                                                                                                                                        .                                                                                      	                                          	                                                                                             -                                                                                                                                                                                                                                  .                                                                                           	                                                                                                                          	-              	                                                                                                                                                                                                                         -                                                                                                                                                                                                                       ,       	                                                                                                                                                                                                                     0                                                                                                                                                                                                                 ,                                                                                                                                                                                                         
                 /                                                                                                                                                                                                                         ,                  	0                                                                                                                                                                                                                                  .                                                                                                                                                                                                                           	    ,                                                                                                                                                                                                                                           -                                                                                                                                                                                                                              #              ,                                                                                                                                                                                                                             0                                                                                                                                                                                                                ,       	                        
  	                                                                                                                                                                                            -                                                                                                                                                                                                           1                             
       ,                                                                                                                                                                                                                              	       ,                                    	 *                                                                                                                                                                                                          /                                                                                                                               
                                                                                    .                                                                                                                                                                                                                               	          -                                                                                                                                                                                                                                  -                                                                                                                                            +	                                                                                                    -                                                                                                                                                                                                                              ,                                                                                                                                                                                                            	                         +        -           !                                                                                                                                                                                                                             -                                                                                                                                                                                                                          ,                                                                                                                                                                                                                     	       ,                                                                                                                                                                                                                                 $                    ,            8                                                                                                                                                                                                                                     /                                                                                                                                                                                                                     -                 
                                                                                                                                                                                                            -                                                                                                                                                                                                                       ,                                                                                                                                                                                                                                       .                                                                                                                                                                                                                            .                                                                                                                                                                                                                                     /                                                                                                                                                                                                                          	      /                                                                                                                                                                                                              0                                                                                                                                                                                                             -                                                                                                                                                                                                                            -                                                                                         	                                                                                                                                 -                                                                                                                                                                                                                                   /                                                                                                                                                                                                        /                                                                                                                                                                                                                	                      -                                                                                                                                                                                                                               -         	    	                                                                                                                                                                                                                     -                                                                                       
                                                                                                                    	         0          	                                                                                                                                                                                                                      ,                                                                                                                                                                                                                               -                                                                                                                                                                                                                            /                                                                                                                                                                                                                0                                                                                                                                                                                                                        	    .                                                                                                                                                                                                                                .                                                                                                                                                                                                                   .                                                                                                                                                                                                                        ,             
                                                                                                                                                                                                              	-                
                                                                                                                                                                                                (                  -               
                                                                                                                                                                                             	            -                                                                                                                          	                                                                                   /      
                                                                                                                                                                                                                              ,                                                                                                                                                                                                                             !               -               $                                                                                                                                                                                                                   -                                                                                        	                                                                                                                              -      	                   
                                                                                                                                                                                             /                                                                                                                                                                                                                      ,                                                                                           	 
                                                                                                                                            /                             	                                                                                                                                                                                                -                                                                                          	                                                                                                                               0                                                                                                                                                                                                        -                                                                                                                                                                                   
                            .                                                                                                                                                                                                                       0                                                                                                                                                                                                                ,                                                                                                                                                                                                                             ,                                  	                                                                                                                                                                                                    .                               
                                                                                                                                                        
                                 -                                                                                                                          	                                                                                           -                                    	                                                                                                                                                                                                  .                                    	                                                                                                                                                                                       /                                                                                                                                                                                                      /    
                	                                                                                                                                                                                                        .         	             	                                                                                                                                                                                           	                 /                                                                                                                                                                                              	                        .                                                                                                                                                                                                                    ,  
                                                                                                                                                                                                                            .                                                                                                                                                                                                                                  .                                                                                                                                
                                                                                            .                                                                                                                                                                                                           
         .                                                                                                                                                                                                                                -                                   	                                                                                                                                                                                              .             	                                                                                                                                                                                                                    0                                                                                                                                                                                                            /           
                                                                                                                                                                                                                            -                                                                                                                             
 
                                                                                         .               	                                                                                                                                                                                         	                       .                                                                                                                                                                                                                  -                                                                                                                                                                                                                 	                     -                                                                                                                                                                                                                                   -                                                                                                                                                                                                                            0                                                                                                                                                                                                                   /                                                                                                                                                                                                                                      -                                                                                                                                                                                                                        	   1                                   	                                                 	                                                                                                                              .                                                                                                                                                                                                                     -     
                                                                                                                                                                                                                            ,                                                                                                                                                                                                                               	      -                                                                                                                                                                                                                        3                                                                                                                                                                                                                    .  	                                                                                                                                                                                                                      .                                                                                                     	                                                                                                                                       ,              !                                                                                                                                                                                                                -                                                                                                                                                                                                                  -                                                                                                                                                                                                                            .                                                                                                                                                                                                                   ,                                    	 	                                                                                                                                                                                                      -                               	                                                          
                                                                                                                                       /                                                                                                                                                                                                                    .                                                                                                                                                                                                            .                                                                                                                                                                                           
                                -   	                                                                                                                           	                                                                                             -                                                                                                                                                                                	                            -                                                                                                                                                                                                                                   "     	   -                                	                                                                                                                                                                                                       /                                	                                                                                                                                                     	                                  ,          
                                                                                                               	                                                                                             ,          
                           	                                                                                                                                                                           	                    
      /                                                                                                                                                                                                                          1                            	                                                                                                                                                                         -                                                                                                                                                                                                                                -                      
                                                                                                                                                                                                              /                                                                                                                                                                                                                        
   -                                                                                                                                                                                                                           -  
                                            
                                                                                                                                                                               /                                                                                                                                                                         	                                0               	                                                                                                                	                                                                                       .                                                                                                                                                                                                                 	-                                                                                                                                    	                                                                                      /                                	 
                                                      
                                                                                                                                      .                                                                                                                                                                                                                          .                                                                                                                                                                                                      	                -                                                                                                                                                                                                                     0                                                                                                                                                                                                   .                                                                                                                                                                                                                                .                                                                                                                                                                                                       
           
    /                                                                                                                                                                                                                /                                                                                                                                                                                                          .                                                                                                                                                                                                                         /                                                                                                                                                                                                               .                                                                                                                                                                                                                          .                                                                                                                                                                                                                 ,                                                                                  
                                                                                                                                      ,                                                                                                                                        
                                                                                          -                                                                                   	                                                                                                                                   .                                                                                                                                                                                                     
      	         ,                                                                                        
                                                                                                                                   .                                                                                                                                                                                                             .        
                                                                                                                                                                                                               -                                                                                    
                                                                                                                            
           -                                                                                                                                                                                                                          1                                                                                                                                                                                                             /                               
                                                                                                                                                                                                  .                                                                                              	                                                                                                                              3                                                                                                                                                                                                           0                               
                                                      
                                                                                                                               .                                                                                                                            
                                                                                   0                                                                                                                                                                                                             	0                                                                                                                                                                                                               0                                                                                                                     	                                                                                      1                                                                                                                                                                                                             /                                                                                                                                                                                                                                	  -                                                                                                                                                                                                                    /                                                                                                                                                                             	                            ,                                                                                                                                                                                                                          .                                                                                                                                                                                                                          	   	    /                                                                                                                                                                                                                  	.                                                                                                                                                                                                          /                                                                                                                                                                                                                          /                                                                                                                                                                                                                 .             
                                                                                                                                                                                                 -                                                                                                                                                                                                                   -                                                                                                                                                                                                                             .                                                                                                                                                                                                  	         -              	                                                                                                                                                                                                         .                                                                                                                                                                                                                         ,                                                                                                                                           
                                                                                    -                                                                                                                                                                                                                         .                                                                                                                                                                                                                          -                                                                                                                                                                                                                 
                  -                                                                                                                                                                                                                              .                                                                                                                                 	                                                                                  -       
     	                                                                                                                                                                                                         .                                                                                                                                                                                                                                   
   .  	           	                                                                                                                                                                                                     2                                                                                                                                                                                                          -                                                                                                                                                                                                                             /                                                                                                                                                                                                                            -  	                               	                                                                                                                                                                                            .                                
                                                                                                                                                                                      .                                                                                     	                                                                                                                                           ,                                                                                                                                                                                                                               .                                                                                    
                                                                                                                                  -                                                                                                                                                                                                                      -                                                                                      
                                                                                                                               .                                                                                                                       	                                                                                      -     
    
     	                                                                                                                                                                                                                     ,                                                                                                                                                                                                               
                       -              	                                                                                                                                                                                                    .                           	                                                                                                                                                                             -                                                                                                                                                                                                                           ,                                                                                                                                                                                                                           1                                                                                                                                                                                                                 -                                                                                                                                                                                                                 0                                                                                                                              
                                                                                   0                                                                                                                                                                                                            0                                                                                                                                                                                                            	1                                                                                                                             
                                                                                         /                                                                                                                                                                                                               .                                                                                                                                                                                                           
                	   .    	            
                                                                                                                                                                                                       1                                                                                                                                                                                                               -                                                                                                                                 
                                                                                              /                                                                                                                                                                                                	                 	   -     	                                                                                                                                                                                                          /         	                    	                                                                                                                                                                            .                                
                                                                                                                                                                                    .                                                                                                                                                                                                           -                                                                                                                                                                                                            -                                                                                                                                                                                                                             -       	                                                                                                                                                                                                        0                                                                                                                                                                                    	                                    ,                                                                                                                                                                                                                       0                                                                                                                                                                                                        .                                                                                                                                                                                                                             ,                                                                                       	                                                                                                                                   -          
                                                                                                                                                                                                                       .                                                                                                                                                                                                             /                                                                                                                                                                                                                      ,                                                                                                                                                                                                                     ,              
                                                                                                                                                                                                              -                                                                                                                                                                                                               	      2       
          	                                                                                                                                                                                               -                                                                                      
                                                                                                                 	                 -                                                                                                                                                                                                                                ,                                                                                                                                                                                                                  
            /    
              	            	                                                                                                                                                                                                    0                                                                                                                                                                                                                       0                                                                                                                                                                                                                       ,                                                                                                                                                                                                                            -                                                                                                                                                                                                                            .                                                                                                                                                                                                                                	    ,                                                                                                                                                                                                           .                                                                                                                                                                                                        ,                                                                                                                                                                                                                              .                                                                                                                                                                                                            
       
           -                                                                                                                                                                                                                       2                                   
                                                                                                                                                                                 -                                                                                                                                                                                                                               -                                                                                           
                                                                                                                                     0                                                                                                                                                                                                                  0                             	                                                    	                                                                                                                                /                                                                                          
                                                                                                                             /                                                                                                                                                                                                     .                                                                                                                                                                                                               /                                                                                                                                                                                                                      .                                                                                                                                                                                        
                       	     -                                                                                                                                                                                                                         -                                                                                                                                                                                                                      0                                                                                                                                                                                                           -                                                                                                                                                                                                                                -                                                                                                                                                                                                                         
   -                                                                                                                                                                                                                   0                                	                                                                                                                                                                               .                                                                                                                                                                                                                         .                                                                                         	                                                                                                              	           /                                                                                                                                                                                                             -                                                                                                                                                                                                                        ,                                                                                                                                                                                                                              2                                                                                                                                                                                                             -            	                                                                                                                                                                                                         .                                                                                                                                                                                                                     
            1                                                                                                                                                                                                                  -                                                                                                                                                                                                                        .                                                                                                                                                                                                                                        .                                                                                                                                                                                                              	          
      0                                                                                                                                                                                                               0                                                                                                                                                                                                             ,         
                                                                                                                                                                                                                   .                                                                                                                                                                                                                                0                                                                                                                                                                                                      	      
.                                                                                                                                                                                                    -                                
                                                                                                                                                                                          ,                                                                                                                                                                                                                 
     $           /         	                                                                                                                                                                                                          .                                                                                                                                                                                                                      .                                                                                                                                                                                                                       -                                                                                                                                                                                          	                               ,                                                                                                                                                                                                       -                                                                                                                                                                                                                  +                   ,                                                                                                                                                                                                                           .                                                                                                                                                                                                                  /                                                                                                                                                                                                                  -                                                                                                                                                                                                                     )     	         -                 !                                                                                                                                                                                                          /                                                                              	                                                                                                                               0     	                                                                                                                                                                                                                  -                                                                                                                                                                                                                       .                                                                                   
                                                                                                                                     .                           	                                                                                                                                                                                         /                                                                                      
                                                                                         	                               1                                                                                                                                                                                              	1                                                                                                                                                                                                            	,                                                                                                                             
                                                                                           .                                                                                                                                                                                                     -                                                                                                                                                                                                                               *     -    
                                                                                                                                                                                                                     /                                                                                                                                                                                 
                                 /                                                                                                                                                                                                                                   /                                                                                                                                                                                                                                   
   ,                                                                                                                                                                                                                             1                                                                                                               	                                                                                         .                                                                                                                                                                                                             0                                                                                                                                                                                                                       
          -                                                                                                                                                                                                                .                                                                                                                                                                                                                              -                                                                                                                                                                                                                                   0                                                                                                                                                                                     
                                 -                                                                                                                                                                                                                 -                                                                                                                                                                                                               .                                                                                                                                                                                                       	                 ,                                                                                                                                                                                                                                        -                                                                                                                                                                                                                                -                                                                                                                                                                                                               .     	                 	                                                                                                                                                                                                                      0                                                                                                                                                                                                                   -                                                                                                                                                                                                                                
    ,                                                                                                                                                                                                               /     	                                                                                                                                                                                                                        	                    0                                                                                                                                                                                                         /                                                                                                                                                                                                                   /                                                                                                                                                                                                            	    .                                                                                                                                                                                                                    1                                                                                                                                                                                                                         ,                                                                                                                                                                                                                      ,                                                                                                                                                                                                               	       .                                                                                                                                                                                                          -                                                                                                                                                                                                                     5                   ,                                                                                                                                                                                                               .                                                                                                                                                                                                                      .                                                                                                                                                                                                               .                                                                                                                                                                                                                          #          	    ,                                                                                                                                                                                                                                  0                                                                                  	                                                                                                             	             .                                                                                                                                                                                                              -                                                                                                                                                                                                              	         	  .                                 	                                                                                                                                                                                        1                                                                                                                                                                                                                        /                                                                                                                                                                                                               -                                                                                                                                                                                                          0                                                                                                                                                                                                       .                                                                                                                                                                                                                 
0                                                                                                                                                                                                          -                                                                                                                                                                                                                         $     /                                                                                                                                                                                                                    .                                                                                                                                                                                                              -                   	                                                                                                              
                                                                                           .                                                                                                                                                                                                                             $           -                                                                                                                                                                                                                       .                                                                                                                                                                                                                  .    	                                                                                                                                                                                                          /                                                                                                                                                                                                                           	           0                                                                                                                                                                                                             -                                                                                       	                                                                                                                                        .                    
                                                                                                                                                                                                              /                                                                                                                                                                                                         .                                                                                                                                                                                                                         .                                                                                                                                                                                                            	   .                	                                                                                                                        	                                                                                          ,                                                                                        
                                                                                                                     	                  -                                                                                                                                                                                                                                        /                                                                                                                                                                                                                  
  /                                                                                                                                                                                                              
    
    .                                                                                                                                                                                                         -                	                                                                                                                                                                                                               ,                                                                                                                                                                                                          
               1                                                                                                                                                                                           	                     0                                                                                                                                                                                                          -                                                                                                                                                                                                                                        /                                                                                                                                                                                                                 2                                                                                                                                                                                                                              -                                                                                                                                                                                                                    /                                                                                       
                                                                                                                               -                                                                                                                                                                                                                       2                                                                                                                                                                                                                /                                                                                                                                                                                                                         7                 /                                                                                                                                                                                                                    0                                                                                                                                                                                                                 0                            	                                                                                                                                                                                    -                                                                                                                                                                                                                        '           -               *                                                                                                                                                                                                                  2                                                                                                                                                                                                              .                                                                                                                                                                                                                  0                                                                                                                                                                                                                     	 1                                                                                           	                                                                                                                                   -                                                                                                                                                                                                                        /                                                                                                                                                                                                            /                                                                                                                                                                                                0                                                                                                                                                                                                              /                                                                                                                                                                                                              -                                                                                                                                                                                                           ,                                                                                                                                                                                                                        "         -                         
                                                                                                                                                                                            	0                                                                                                                                                                                                        ,               	                                                                                                                                                                                                       -                                                                                                                                                                                                                                     .                                                                                                                                                                                                                         ,                                                                                                                                                                                                              0                                                                                                                                                                                                             -                     	                                                                                                                                                                                     	       	       	           0                                                                                                                                 
                                                                         .            	                                                                                                                                                                                                                ,                                            	                                                                                                                                                                                    